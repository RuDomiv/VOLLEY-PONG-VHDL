LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

PACKAGE ImagePackage IS
    
	 TYPE ImageMatrix IS ARRAY (NATURAL RANGE <>, NATURAL RANGE <>) OF STD_logic_vector(7 DOWNTO 0);
	 
	 CONSTANT pokeR : ImageMatrix(0 TO 39, 0 TO 39) := (
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" ),
( x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" ),
( x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" ),
( x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"00" , x"00" , x"00" , x"00" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" ),
( x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" ),
( x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" ),
( x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" )
);


CONSTANT pokeG : ImageMatrix(0 TO 39, 0 TO 39) := (
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" ),
( x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" ),
( x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" ),
( x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"00" , x"00" , x"00" , x"00" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" ),
( x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" ),
( x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" ),
( x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" )
);



CONSTANT pokeB : ImageMatrix(0 TO 39, 0 TO 39) := (
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" ),
( x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" ),
( x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" ),
( x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" ),
( x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"00" , x"00" , x"00" , x"00" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" ),
( x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" ),
( x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" ),
( x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" ),
( x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" )
);


-- Player 1 ASSETS
-----------------------------------------------------------------------------------------------------------------------------------------------

CONSTANT Player1R : ImageMatrix(0 TO 24, 0 TO 99) := (
( x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" ),
( x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" ),
( x"3F" , x"3F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"3F" , x"3F" ),
( x"3F" , x"3F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"02" , x"03" , x"03" , x"03" , x"03" , x"03" , x"02" , x"01" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"01" , x"02" , x"02" , x"01" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"3F" , x"3F" ),
( x"3F" , x"3F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"05" , x"22" , x"34" , x"34" , x"34" , x"34" , x"34" , x"2E" , x"23" , x"11" , x"02" , x"00" , x"00" , x"00" , x"00" , x"00" , x"01" , x"08" , x"1C" , x"2E" , x"2F" , x"10" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"3F" , x"3F" ),
( x"3F" , x"3F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"09" , x"2C" , x"3F" , x"36" , x"2F" , x"2E" , x"31" , x"36" , x"3B" , x"33" , x"17" , x"03" , x"00" , x"00" , x"00" , x"06" , x"16" , x"2B" , x"39" , x"3E" , x"3A" , x"14" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"3F" , x"3F" ),
( x"3F" , x"3F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"09" , x"2D" , x"3F" , x"27" , x"0E" , x"0B" , x"0C" , x"16" , x"30" , x"3D" , x"35" , x"0D" , x"01" , x"00" , x"01" , x"21" , x"36" , x"39" , x"2C" , x"3B" , x"3A" , x"15" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"3F" , x"3F" ),
( x"3F" , x"3F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"09" , x"2D" , x"3F" , x"23" , x"04" , x"00" , x"00" , x"01" , x"17" , x"36" , x"3E" , x"1B" , x"03" , x"00" , x"02" , x"2E" , x"2B" , x"15" , x"09" , x"35" , x"3A" , x"15" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"3F" , x"3F" ),
( x"3F" , x"3F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"09" , x"2D" , x"3F" , x"23" , x"04" , x"00" , x"00" , x"00" , x"0C" , x"30" , x"3E" , x"22" , x"04" , x"00" , x"01" , x"0D" , x"08" , x"02" , x"02" , x"34" , x"3A" , x"15" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"3F" , x"3F" ),
( x"3F" , x"3F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"09" , x"2D" , x"3F" , x"23" , x"04" , x"00" , x"00" , x"00" , x"0C" , x"30" , x"3E" , x"22" , x"04" , x"00" , x"00" , x"01" , x"00" , x"00" , x"02" , x"34" , x"3A" , x"15" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"3F" , x"3F" ),
( x"3F" , x"3F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"09" , x"2D" , x"3F" , x"23" , x"04" , x"00" , x"00" , x"00" , x"13" , x"36" , x"3E" , x"1B" , x"03" , x"00" , x"00" , x"00" , x"00" , x"00" , x"02" , x"34" , x"3A" , x"15" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"3F" , x"3F" ),
( x"3F" , x"3F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"09" , x"2D" , x"3F" , x"24" , x"06" , x"02" , x"03" , x"0A" , x"28" , x"3C" , x"36" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"02" , x"34" , x"3A" , x"15" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"3F" , x"3F" ),
( x"3F" , x"3F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"09" , x"2D" , x"3F" , x"30" , x"21" , x"1F" , x"22" , x"2F" , x"3A" , x"36" , x"1A" , x"03" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"02" , x"34" , x"3A" , x"15" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"3F" , x"3F" ),
( x"3F" , x"3F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"09" , x"2D" , x"3F" , x"3D" , x"3B" , x"3B" , x"3B" , x"37" , x"2C" , x"18" , x"05" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"02" , x"34" , x"3A" , x"15" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"3F" , x"3F" ),
( x"3F" , x"3F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"09" , x"2D" , x"3F" , x"2D" , x"18" , x"15" , x"14" , x"10" , x"09" , x"03" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"02" , x"34" , x"3A" , x"15" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"3F" , x"3F" ),
( x"3F" , x"3F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"09" , x"2D" , x"3F" , x"23" , x"04" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"02" , x"34" , x"3A" , x"15" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"3F" , x"3F" ),
( x"3F" , x"3F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"09" , x"2D" , x"3F" , x"23" , x"04" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"02" , x"34" , x"3A" , x"15" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"3F" , x"3F" ),
( x"3F" , x"3F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"09" , x"2D" , x"3F" , x"23" , x"04" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"02" , x"34" , x"3A" , x"15" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"3F" , x"3F" ),
( x"3F" , x"3F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"09" , x"2D" , x"3F" , x"23" , x"04" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"09" , x"10" , x"10" , x"12" , x"37" , x"3A" , x"1F" , x"10" , x"10" , x"09" , x"01" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"3F" , x"3F" ),
( x"3F" , x"3F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"09" , x"2C" , x"3F" , x"23" , x"04" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"01" , x"26" , x"35" , x"37" , x"37" , x"3E" , x"3E" , x"39" , x"37" , x"37" , x"26" , x"08" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"3F" , x"3F" ),
( x"3F" , x"3F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"05" , x"1D" , x"2B" , x"16" , x"03" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"01" , x"1D" , x"2A" , x"2B" , x"2B" , x"2B" , x"2B" , x"2B" , x"2B" , x"2B" , x"1D" , x"06" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"3F" , x"3F" ),
( x"3F" , x"3F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"01" , x"03" , x"05" , x"02" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"03" , x"05" , x"05" , x"05" , x"05" , x"05" , x"05" , x"05" , x"05" , x"03" , x"01" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"3F" , x"3F" ),
( x"3F" , x"3F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"3F" , x"3F" ),
( x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" ),
( x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" , x"3F" )
);

CONSTANT Player1G : ImageMatrix(0 TO 24, 0 TO 99) := (
( x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" ),
( x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" ),
( x"48" , x"48" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"48" , x"48" ),
( x"48" , x"48" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A1" , x"A0" , x"9E" , x"9E" , x"9E" , x"9E" , x"9E" , x"9F" , x"A0" , x"A1" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A0" , x"9F" , x"9F" , x"A1" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"48" , x"48" ),
( x"48" , x"48" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"9A" , x"71" , x"58" , x"58" , x"58" , x"58" , x"58" , x"60" , x"70" , x"8B" , x"9F" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A0" , x"96" , x"7A" , x"60" , x"60" , x"8B" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"48" , x"48" ),
( x"48" , x"48" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"96" , x"63" , x"49" , x"55" , x"5F" , x"60" , x"5D" , x"54" , x"4D" , x"58" , x"82" , x"9D" , x"A2" , x"A2" , x"A2" , x"9A" , x"82" , x"65" , x"50" , x"4A" , x"50" , x"85" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"48" , x"48" ),
( x"48" , x"48" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"95" , x"62" , x"49" , x"6B" , x"8D" , x"93" , x"90" , x"82" , x"5E" , x"4A" , x"56" , x"91" , x"A1" , x"A2" , x"A0" , x"72" , x"56" , x"52" , x"63" , x"4E" , x"4F" , x"84" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"48" , x"48" ),
( x"48" , x"48" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"95" , x"62" , x"49" , x"70" , x"9C" , x"A2" , x"A2" , x"A0" , x"83" , x"54" , x"49" , x"7A" , x"9D" , x"A2" , x"A0" , x"60" , x"64" , x"85" , x"95" , x"57" , x"4F" , x"84" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"48" , x"48" ),
( x"48" , x"48" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"95" , x"62" , x"49" , x"70" , x"9C" , x"A2" , x"A2" , x"A2" , x"90" , x"5D" , x"48" , x"72" , x"9C" , x"A2" , x"A2" , x"8F" , x"97" , x"A0" , x"9F" , x"58" , x"4F" , x"84" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"48" , x"48" ),
( x"48" , x"48" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"95" , x"62" , x"49" , x"70" , x"9C" , x"A2" , x"A2" , x"A2" , x"91" , x"5E" , x"48" , x"71" , x"9C" , x"A2" , x"A2" , x"A0" , x"A1" , x"A2" , x"9F" , x"58" , x"4F" , x"84" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"48" , x"48" ),
( x"48" , x"48" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"95" , x"62" , x"49" , x"70" , x"9C" , x"A2" , x"A2" , x"A2" , x"88" , x"55" , x"49" , x"7B" , x"9E" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"9F" , x"58" , x"4F" , x"84" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"48" , x"48" ),
( x"48" , x"48" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"95" , x"62" , x"49" , x"70" , x"99" , x"9F" , x"9F" , x"94" , x"68" , x"4B" , x"55" , x"91" , x"A1" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"9F" , x"58" , x"4F" , x"84" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"48" , x"48" ),
( x"48" , x"48" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"95" , x"62" , x"48" , x"5D" , x"73" , x"76" , x"71" , x"5F" , x"4F" , x"55" , x"7D" , x"9D" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"9F" , x"58" , x"4F" , x"84" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"48" , x"48" ),
( x"48" , x"48" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"95" , x"62" , x"48" , x"4A" , x"4D" , x"4E" , x"4E" , x"53" , x"64" , x"81" , x"9B" , x"A1" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"9F" , x"58" , x"4F" , x"84" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"48" , x"48" ),
( x"48" , x"48" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"95" , x"62" , x"49" , x"63" , x"80" , x"83" , x"85" , x"8A" , x"94" , x"9F" , x"A1" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"9F" , x"58" , x"4F" , x"84" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"48" , x"48" ),
( x"48" , x"48" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"95" , x"62" , x"49" , x"70" , x"9C" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"9F" , x"58" , x"4F" , x"84" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"48" , x"48" ),
( x"48" , x"48" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"95" , x"62" , x"49" , x"70" , x"9C" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"9F" , x"58" , x"4F" , x"84" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"48" , x"48" ),
( x"48" , x"48" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"95" , x"62" , x"49" , x"70" , x"9C" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"9F" , x"58" , x"4F" , x"84" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"48" , x"48" ),
( x"48" , x"48" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"95" , x"62" , x"49" , x"70" , x"9C" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A1" , x"95" , x"8B" , x"8A" , x"88" , x"54" , x"4E" , x"76" , x"8A" , x"8A" , x"95" , x"A1" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"48" , x"48" ),
( x"48" , x"48" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"95" , x"63" , x"49" , x"70" , x"9C" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A1" , x"6C" , x"55" , x"54" , x"53" , x"4A" , x"49" , x"51" , x"54" , x"54" , x"6C" , x"97" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"48" , x"48" ),
( x"48" , x"48" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"9B" , x"78" , x"65" , x"82" , x"9D" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A0" , x"78" , x"67" , x"65" , x"65" , x"65" , x"65" , x"65" , x"65" , x"65" , x"78" , x"9A" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"48" , x"48" ),
( x"48" , x"48" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"9D" , x"9B" , x"9F" , x"A1" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"9D" , x"9B" , x"9B" , x"9B" , x"9B" , x"9B" , x"9B" , x"9B" , x"9B" , x"9D" , x"A1" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"48" , x"48" ),
( x"48" , x"48" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"48" , x"48" ),
( x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" ),
( x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" , x"48" )
);

CONSTANT Player1B : ImageMatrix(0 TO 24, 0 TO 99) := (
( x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" ),
( x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" ),
( x"CC" , x"CC" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CC" , x"CC" ),
( x"CC" , x"CC" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"E7" , x"E7" , x"E7" , x"E7" , x"E7" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"E7" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CC" , x"CC" ),
( x"CC" , x"CC" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"D8" , x"D1" , x"D1" , x"D1" , x"D1" , x"D1" , x"D4" , x"D9" , x"E1" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E4" , x"DC" , x"D3" , x"D3" , x"E1" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CC" , x"CC" ),
( x"CC" , x"CC" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E4" , x"D4" , x"CC" , x"D0" , x"D3" , x"D4" , x"D3" , x"CF" , x"CE" , x"D1" , x"DD" , x"E6" , x"E8" , x"E8" , x"E8" , x"E5" , x"DE" , x"D6" , x"CE" , x"CD" , x"CE" , x"DF" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CC" , x"CC" ),
( x"CC" , x"CC" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E3" , x"D3" , x"CC" , x"D7" , x"E1" , x"E3" , x"E3" , x"DE" , x"D2" , x"CD" , x"D0" , x"E3" , x"E7" , x"E8" , x"E7" , x"D9" , x"D0" , x"D0" , x"D4" , x"CD" , x"CE" , x"DE" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CC" , x"CC" ),
( x"CC" , x"CC" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E3" , x"D3" , x"CC" , x"DA" , x"E7" , x"E8" , x"E8" , x"E8" , x"DE" , x"D0" , x"CC" , x"DC" , x"E7" , x"E8" , x"E8" , x"D3" , x"D5" , x"DF" , x"E4" , x"D1" , x"CE" , x"DE" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CC" , x"CC" ),
( x"CC" , x"CC" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E3" , x"D3" , x"CC" , x"DA" , x"E7" , x"E8" , x"E8" , x"E8" , x"E3" , x"D3" , x"CC" , x"D9" , x"E7" , x"E8" , x"E8" , x"E2" , x"E5" , x"E8" , x"E7" , x"D2" , x"CE" , x"DE" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CC" , x"CC" ),
( x"CC" , x"CC" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E3" , x"D3" , x"CC" , x"DA" , x"E7" , x"E8" , x"E8" , x"E8" , x"E2" , x"D2" , x"CC" , x"D9" , x"E6" , x"E8" , x"E8" , x"E7" , x"E8" , x"E8" , x"E7" , x"D2" , x"CE" , x"DE" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CC" , x"CC" ),
( x"CC" , x"CC" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E3" , x"D3" , x"CC" , x"DA" , x"E7" , x"E8" , x"E8" , x"E8" , x"E0" , x"CF" , x"CC" , x"DC" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"D2" , x"CE" , x"DE" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CC" , x"CC" ),
( x"CC" , x"CC" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E3" , x"D3" , x"CC" , x"D9" , x"E5" , x"E8" , x"E7" , x"E4" , x"D6" , x"CC" , x"D0" , x"E2" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"D2" , x"CE" , x"DE" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CC" , x"CC" ),
( x"CC" , x"CC" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E3" , x"D3" , x"CC" , x"D2" , x"D9" , x"D9" , x"DA" , x"D3" , x"CE" , x"D1" , x"DD" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"D2" , x"CE" , x"DE" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CC" , x"CC" ),
( x"CC" , x"CC" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E3" , x"D3" , x"CC" , x"CC" , x"CE" , x"CE" , x"CE" , x"CF" , x"D5" , x"DE" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"D2" , x"CE" , x"DE" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CC" , x"CC" ),
( x"CC" , x"CC" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E3" , x"D3" , x"CD" , x"D4" , x"DD" , x"DE" , x"DF" , x"E1" , x"E3" , x"E7" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"D2" , x"CE" , x"DE" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CC" , x"CC" ),
( x"CC" , x"CC" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E3" , x"D3" , x"CC" , x"DA" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"D2" , x"CE" , x"DE" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CC" , x"CC" ),
( x"CC" , x"CC" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E3" , x"D3" , x"CC" , x"DA" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"D2" , x"CE" , x"DE" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CC" , x"CC" ),
( x"CC" , x"CC" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E3" , x"D3" , x"CC" , x"DA" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"D2" , x"CE" , x"DE" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CC" , x"CC" ),
( x"CC" , x"CC" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E3" , x"D3" , x"CC" , x"DA" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E4" , x"E1" , x"E0" , x"E0" , x"D0" , x"CD" , x"DA" , x"E0" , x"E0" , x"E4" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CC" , x"CC" ),
( x"CC" , x"CC" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E4" , x"D4" , x"CC" , x"DA" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"D8" , x"D0" , x"CF" , x"D0" , x"CC" , x"CC" , x"CF" , x"CF" , x"CF" , x"D8" , x"E5" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CC" , x"CC" ),
( x"CC" , x"CC" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"DC" , x"D5" , x"DE" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"DB" , x"D6" , x"D5" , x"D5" , x"D5" , x"D5" , x"D5" , x"D5" , x"D5" , x"DB" , x"E5" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CC" , x"CC" ),
( x"CC" , x"CC" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"E6" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"E6" , x"E6" , x"E6" , x"E6" , x"E6" , x"E6" , x"E6" , x"E6" , x"E6" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CC" , x"CC" ),
( x"CC" , x"CC" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CC" , x"CC" ),
( x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" ),
( x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" , x"CC" )
);






-- player 2 assETS
-----------------------------------------------------------------------------------------------------------------------------------------------

CONSTANT Player2R : ImageMatrix(0 TO 24, 0 TO 99) := (
( x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" ),
( x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" ),
( x"88" , x"88" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"88" , x"88" ),
( x"88" , x"88" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"EC" , x"E9" , x"E9" , x"E9" , x"E9" , x"E9" , x"E9" , x"EA" , x"EB" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"EC" , x"EB" , x"EA" , x"EA" , x"E9" , x"EA" , x"EB" , x"EC" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"88" , x"88" ),
( x"88" , x"88" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"E6" , x"B9" , x"9A" , x"9A" , x"9A" , x"9A" , x"99" , x"A4" , x"B9" , x"D4" , x"EA" , x"ED" , x"ED" , x"ED" , x"EA" , x"D9" , x"BE" , x"AA" , x"9C" , x"9A" , x"A3" , x"B9" , x"D9" , x"EA" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"88" , x"88" ),
( x"88" , x"88" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"E3" , x"AA" , x"88" , x"97" , x"A5" , x"A7" , x"A3" , x"98" , x"91" , x"9E" , x"CC" , x"E9" , x"ED" , x"ED" , x"D8" , x"A5" , x"92" , x"98" , x"9C" , x"97" , x"8D" , x"8E" , x"A2" , x"D5" , x"EB" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"88" , x"88" ),
( x"88" , x"88" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"E2" , x"A9" , x"89" , x"B4" , x"D9" , x"DF" , x"DC" , x"CE" , x"A3" , x"8B" , x"9A" , x"DA" , x"EC" , x"ED" , x"C8" , x"A6" , x"BB" , x"D0" , x"D6" , x"D2" , x"B1" , x"8F" , x"8B" , x"B2" , x"E5" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"88" , x"88" ),
( x"88" , x"88" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"E2" , x"A9" , x"88" , x"BA" , x"E6" , x"ED" , x"ED" , x"EA" , x"CD" , x"98" , x"8A" , x"C6" , x"E9" , x"ED" , x"E4" , x"DF" , x"E8" , x"EC" , x"ED" , x"ED" , x"DF" , x"A5" , x"88" , x"9E" , x"DC" , x"EC" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"88" , x"88" ),
( x"88" , x"88" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"E2" , x"A9" , x"88" , x"BA" , x"E6" , x"ED" , x"ED" , x"ED" , x"DD" , x"A4" , x"89" , x"BC" , x"E7" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"EB" , x"AF" , x"88" , x"9B" , x"D7" , x"EC" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"88" , x"88" ),
( x"88" , x"88" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"E2" , x"A9" , x"88" , x"BA" , x"E6" , x"ED" , x"ED" , x"ED" , x"DD" , x"A3" , x"89" , x"BB" , x"E7" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"EA" , x"AD" , x"88" , x"9F" , x"DD" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"88" , x"88" ),
( x"88" , x"88" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"E2" , x"A9" , x"88" , x"BA" , x"E6" , x"ED" , x"ED" , x"ED" , x"D0" , x"99" , x"8A" , x"C7" , x"E9" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"DF" , x"A3" , x"89" , x"AF" , x"E4" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"88" , x"88" ),
( x"88" , x"88" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"E2" , x"A9" , x"88" , x"B8" , x"E4" , x"EA" , x"EA" , x"DE" , x"B0" , x"8C" , x"99" , x"DB" , x"EC" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"E9" , x"C4" , x"92" , x"8E" , x"C9" , x"EA" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"88" , x"88" ),
( x"88" , x"88" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"E2" , x"A9" , x"89" , x"A5" , x"BE" , x"C0" , x"BC" , x"A5" , x"90" , x"98" , x"C8" , x"E8" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"DA" , x"A5" , x"8C" , x"B2" , x"E1" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"88" , x"88" ),
( x"88" , x"88" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"E2" , x"A9" , x"88" , x"8B" , x"8F" , x"8F" , x"91" , x"98" , x"AB" , x"CB" , x"E6" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"E3" , x"B1" , x"90" , x"A2" , x"D8" , x"EB" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"88" , x"88" ),
( x"88" , x"88" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"E2" , x"A9" , x"89" , x"AA" , x"C7" , x"CB" , x"CC" , x"D4" , x"E0" , x"EA" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"E5" , x"B2" , x"8F" , x"9C" , x"D0" , x"E9" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"88" , x"88" ),
( x"88" , x"88" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"E2" , x"A9" , x"88" , x"BA" , x"E6" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"EC" , x"E3" , x"B3" , x"8D" , x"97" , x"C9" , x"E8" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"88" , x"88" ),
( x"88" , x"88" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"E2" , x"A9" , x"88" , x"BA" , x"E6" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"E4" , x"BD" , x"93" , x"97" , x"C7" , x"E6" , x"EC" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"88" , x"88" ),
( x"88" , x"88" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"E2" , x"A9" , x"88" , x"BA" , x"E6" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"E8" , x"BE" , x"95" , x"9B" , x"C9" , x"E7" , x"EC" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"88" , x"88" ),
( x"88" , x"88" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"E2" , x"A9" , x"88" , x"BA" , x"E6" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"C5" , x"96" , x"8E" , x"AC" , x"C5" , x"C9" , x"C9" , x"C9" , x"C9" , x"CA" , x"DA" , x"EB" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"88" , x"88" ),
( x"88" , x"88" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"E3" , x"A9" , x"88" , x"BA" , x"E6" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"A7" , x"8A" , x"8A" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"B3" , x"E5" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"88" , x"88" ),
( x"88" , x"88" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"E7" , x"BF" , x"A9" , x"CD" , x"E9" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"C3" , x"AB" , x"A8" , x"A8" , x"A8" , x"A8" , x"A8" , x"A8" , x"A8" , x"A9" , x"C6" , x"E9" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"88" , x"88" ),
( x"88" , x"88" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"EC" , x"E8" , x"E5" , x"EA" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"E8" , x"E5" , x"E5" , x"E5" , x"E5" , x"E5" , x"E5" , x"E5" , x"E5" , x"E4" , x"E9" , x"EC" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"88" , x"88" ),
( x"88" , x"88" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"88" , x"88" ),
( x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" ),
( x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" , x"88" )
);

CONSTANT Player2G : ImageMatrix(0 TO 24, 0 TO 99) := (
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"00" , x"00" ),
( x"00" , x"00" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1B" , x"1B" , x"1B" , x"1B" , x"1B" , x"1B" , x"1B" , x"1B" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1B" , x"1B" , x"1B" , x"1B" , x"1B" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"00" , x"00" ),
( x"00" , x"00" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1A" , x"0E" , x"05" , x"05" , x"05" , x"05" , x"05" , x"08" , x"0E" , x"15" , x"1B" , x"1C" , x"1C" , x"1C" , x"1B" , x"16" , x"0F" , x"09" , x"06" , x"05" , x"07" , x"0E" , x"16" , x"1B" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"00" , x"00" ),
( x"00" , x"00" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"19" , x"09" , x"00" , x"04" , x"08" , x"09" , x"07" , x"05" , x"02" , x"06" , x"13" , x"1B" , x"1C" , x"1C" , x"16" , x"08" , x"03" , x"05" , x"06" , x"04" , x"01" , x"02" , x"07" , x"15" , x"1B" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"00" , x"00" ),
( x"00" , x"00" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"19" , x"09" , x"00" , x"0C" , x"17" , x"18" , x"17" , x"13" , x"08" , x"01" , x"05" , x"17" , x"1C" , x"1C" , x"12" , x"08" , x"0E" , x"14" , x"16" , x"14" , x"0B" , x"02" , x"01" , x"0C" , x"1A" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"00" , x"00" ),
( x"00" , x"00" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"19" , x"09" , x"00" , x"0E" , x"1A" , x"1C" , x"1C" , x"1B" , x"13" , x"05" , x"00" , x"11" , x"1B" , x"1C" , x"1A" , x"18" , x"1B" , x"1C" , x"1C" , x"1C" , x"18" , x"08" , x"00" , x"06" , x"17" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"00" , x"00" ),
( x"00" , x"00" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"19" , x"09" , x"00" , x"0E" , x"1A" , x"1C" , x"1C" , x"1C" , x"17" , x"08" , x"00" , x"0E" , x"1A" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"0B" , x"00" , x"05" , x"16" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"00" , x"00" ),
( x"00" , x"00" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"19" , x"09" , x"00" , x"0E" , x"1A" , x"1C" , x"1C" , x"1C" , x"17" , x"08" , x"00" , x"0E" , x"1A" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1B" , x"0A" , x"00" , x"06" , x"18" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"00" , x"00" ),
( x"00" , x"00" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"19" , x"09" , x"00" , x"0E" , x"1A" , x"1C" , x"1C" , x"1C" , x"14" , x"05" , x"00" , x"11" , x"1B" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"18" , x"08" , x"00" , x"0B" , x"1A" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"00" , x"00" ),
( x"00" , x"00" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"19" , x"09" , x"00" , x"0E" , x"1A" , x"1B" , x"1B" , x"18" , x"0B" , x"01" , x"05" , x"17" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1B" , x"11" , x"03" , x"02" , x"12" , x"1B" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"00" , x"00" ),
( x"00" , x"00" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"19" , x"09" , x"00" , x"08" , x"0F" , x"10" , x"0E" , x"08" , x"02" , x"05" , x"12" , x"1B" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"17" , x"08" , x"01" , x"0B" , x"19" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"00" , x"00" ),
( x"00" , x"00" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"19" , x"09" , x"00" , x"01" , x"02" , x"02" , x"02" , x"05" , x"0A" , x"13" , x"1A" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"19" , x"0B" , x"02" , x"07" , x"16" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"00" , x"00" ),
( x"00" , x"00" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"19" , x"09" , x"00" , x"09" , x"11" , x"13" , x"13" , x"15" , x"18" , x"1B" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"19" , x"0C" , x"02" , x"06" , x"14" , x"1B" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"00" , x"00" ),
( x"00" , x"00" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"19" , x"09" , x"00" , x"0E" , x"1A" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"19" , x"0C" , x"02" , x"04" , x"12" , x"1B" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"00" , x"00" ),
( x"00" , x"00" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"19" , x"09" , x"00" , x"0E" , x"1A" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1A" , x"0F" , x"03" , x"04" , x"11" , x"1A" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"00" , x"00" ),
( x"00" , x"00" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"19" , x"09" , x"00" , x"0E" , x"1A" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1B" , x"0F" , x"04" , x"05" , x"12" , x"1A" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"00" , x"00" ),
( x"00" , x"00" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"19" , x"09" , x"00" , x"0E" , x"1A" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"11" , x"04" , x"02" , x"0A" , x"11" , x"12" , x"12" , x"12" , x"12" , x"12" , x"17" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"00" , x"00" ),
( x"00" , x"00" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"19" , x"09" , x"00" , x"0E" , x"1A" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"09" , x"00" , x"00" , x"02" , x"03" , x"03" , x"03" , x"03" , x"03" , x"03" , x"0C" , x"19" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"00" , x"00" ),
( x"00" , x"00" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1A" , x"0F" , x"09" , x"13" , x"1B" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"10" , x"0A" , x"09" , x"09" , x"09" , x"09" , x"09" , x"09" , x"09" , x"09" , x"11" , x"1B" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"00" , x"00" ),
( x"00" , x"00" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1B" , x"1A" , x"1B" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1B" , x"1A" , x"1A" , x"1A" , x"1A" , x"1A" , x"1A" , x"1A" , x"1A" , x"1A" , x"1B" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"00" , x"00" ),
( x"00" , x"00" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" )
);

CONSTANT Player2B : ImageMatrix(0 TO 24, 0 TO 99) := (
( x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" ),
( x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" ),
( x"15" , x"15" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"15" , x"15" ),
( x"15" , x"15" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"23" , x"23" , x"23" , x"23" , x"23" , x"24" , x"23" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"23" , x"24" , x"24" , x"23" , x"24" , x"23" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"15" , x"15" ),
( x"15" , x"15" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"23" , x"1D" , x"18" , x"18" , x"18" , x"18" , x"18" , x"19" , x"1D" , x"21" , x"24" , x"24" , x"24" , x"24" , x"23" , x"21" , x"1D" , x"1A" , x"18" , x"17" , x"1A" , x"1D" , x"21" , x"23" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"15" , x"15" ),
( x"15" , x"15" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"22" , x"1A" , x"15" , x"18" , x"19" , x"1A" , x"19" , x"17" , x"16" , x"18" , x"1F" , x"24" , x"24" , x"24" , x"20" , x"19" , x"17" , x"18" , x"18" , x"18" , x"16" , x"16" , x"19" , x"20" , x"23" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"15" , x"15" ),
( x"15" , x"15" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"23" , x"1A" , x"15" , x"1C" , x"21" , x"22" , x"22" , x"20" , x"19" , x"15" , x"17" , x"22" , x"24" , x"24" , x"1E" , x"1A" , x"1D" , x"20" , x"21" , x"20" , x"1C" , x"15" , x"16" , x"1B" , x"23" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"15" , x"15" ),
( x"15" , x"15" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"23" , x"1A" , x"15" , x"1C" , x"23" , x"24" , x"24" , x"23" , x"20" , x"18" , x"16" , x"1E" , x"24" , x"24" , x"23" , x"22" , x"23" , x"24" , x"24" , x"24" , x"22" , x"19" , x"15" , x"19" , x"22" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"15" , x"15" ),
( x"15" , x"15" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"23" , x"1A" , x"15" , x"1C" , x"23" , x"24" , x"24" , x"24" , x"21" , x"19" , x"15" , x"1D" , x"23" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"1B" , x"15" , x"17" , x"20" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"15" , x"15" ),
( x"15" , x"15" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"23" , x"1A" , x"15" , x"1C" , x"23" , x"24" , x"24" , x"24" , x"21" , x"19" , x"15" , x"1C" , x"23" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"1A" , x"15" , x"18" , x"21" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"15" , x"15" ),
( x"15" , x"15" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"23" , x"1A" , x"15" , x"1C" , x"23" , x"24" , x"24" , x"24" , x"20" , x"18" , x"16" , x"1E" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"22" , x"19" , x"15" , x"1B" , x"23" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"15" , x"15" ),
( x"15" , x"15" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"23" , x"1A" , x"15" , x"1D" , x"23" , x"24" , x"24" , x"22" , x"1B" , x"16" , x"18" , x"21" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"1D" , x"17" , x"16" , x"1F" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"15" , x"15" ),
( x"15" , x"15" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"23" , x"1A" , x"15" , x"19" , x"1D" , x"1D" , x"1D" , x"19" , x"16" , x"17" , x"1F" , x"23" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"21" , x"19" , x"16" , x"1B" , x"22" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"15" , x"15" ),
( x"15" , x"15" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"23" , x"1A" , x"15" , x"15" , x"16" , x"16" , x"16" , x"18" , x"1A" , x"1F" , x"23" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"22" , x"1B" , x"16" , x"18" , x"21" , x"23" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"15" , x"15" ),
( x"15" , x"15" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"23" , x"1A" , x"15" , x"1A" , x"1E" , x"1F" , x"1F" , x"20" , x"22" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"23" , x"1B" , x"16" , x"17" , x"20" , x"23" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"15" , x"15" ),
( x"15" , x"15" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"23" , x"1A" , x"15" , x"1C" , x"23" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"22" , x"1C" , x"15" , x"18" , x"1F" , x"23" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"15" , x"15" ),
( x"15" , x"15" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"23" , x"1A" , x"15" , x"1C" , x"23" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"23" , x"1D" , x"17" , x"18" , x"1E" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"15" , x"15" ),
( x"15" , x"15" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"23" , x"1A" , x"15" , x"1C" , x"23" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"23" , x"1C" , x"17" , x"18" , x"1E" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"15" , x"15" ),
( x"15" , x"15" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"23" , x"1A" , x"15" , x"1C" , x"23" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"1F" , x"17" , x"16" , x"1B" , x"1F" , x"1E" , x"1E" , x"1E" , x"1E" , x"1F" , x"21" , x"23" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"15" , x"15" ),
( x"15" , x"15" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"22" , x"1A" , x"15" , x"1C" , x"23" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"1A" , x"16" , x"16" , x"17" , x"17" , x"17" , x"17" , x"17" , x"17" , x"16" , x"1B" , x"23" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"15" , x"15" ),
( x"15" , x"15" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"23" , x"1D" , x"1A" , x"1F" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"1E" , x"1A" , x"1A" , x"1A" , x"1A" , x"1A" , x"1A" , x"1A" , x"1A" , x"1A" , x"1E" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"15" , x"15" ),
( x"15" , x"15" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"23" , x"23" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"23" , x"23" , x"23" , x"23" , x"23" , x"23" , x"23" , x"23" , x"23" , x"23" , x"23" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"15" , x"15" ),
( x"15" , x"15" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"15" , x"15" ),
( x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" ),
( x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" , x"15" )
);



-- Net ASSETS
--------------------------------------------------------------------------------------------------------------------------------------------------
CONSTANT NetR : ImageMatrix(0 TO 299, 0 TO 29) := (
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" )
);

CONSTANT NetG : ImageMatrix(0 TO 299, 0 TO 29) := (
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" )
);

CONSTANT NetB : ImageMatrix(0 TO 299, 0 TO 29) := (
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" )
);


-- Separator
----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------

CONSTANT SEPARATORR : ImageMatrix(0 TO 9, 0 TO 799) := (
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" )
);

CONSTANT SEPARATORG : ImageMatrix(0 TO 9, 0 TO 799) := (
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" )
);

CONSTANT SEPARATORB : ImageMatrix(0 TO 9, 0 TO 799) := (
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" )
);

-- Numeros
----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------

--Numero 0
CONSTANT R0 : ImageMatrix(0 TO 39, 0 TO 29) := (
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" )
);

CONSTANT G0 : ImageMatrix(0 TO 39, 0 TO 29) := (
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" )
);

CONSTANT B0 : ImageMatrix(0 TO 39, 0 TO 29) := (
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" )
);

--Numero 1

CONSTANT R1 : ImageMatrix(0 TO 39, 0 TO 29) := (
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" )
);

CONSTANT G1 : ImageMatrix(0 TO 39, 0 TO 29) := (
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" )
);

CONSTANT B1 : ImageMatrix(0 TO 39, 0 TO 29) := (
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" )
);


--Numero 2

CONSTANT R2 : ImageMatrix(0 TO 39, 0 TO 29) := (
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" )
);

CONSTANT G2 : ImageMatrix(0 TO 39, 0 TO 29) := (
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" )
);

CONSTANT B2 : ImageMatrix(0 TO 39, 0 TO 29) := (
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" )
);



--Numero 3

CONSTANT R3 : ImageMatrix(0 TO 39, 0 TO 29) := (
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" )
);

CONSTANT G3 : ImageMatrix(0 TO 39, 0 TO 29) := (
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" )
);

CONSTANT B3 : ImageMatrix(0 TO 39, 0 TO 29) := (
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" )
);

--Numero 4
CONSTANT R4 : ImageMatrix(0 TO 39, 0 TO 29) := (
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" )
);

CONSTANT G4 : ImageMatrix(0 TO 39, 0 TO 29) := (
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" )
);

CONSTANT B4 : ImageMatrix(0 TO 39, 0 TO 29) := (
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" )
);

--Numero 5

CONSTANT R5 : ImageMatrix(0 TO 39, 0 TO 29) := (
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" )
);

CONSTANT G5 : ImageMatrix(0 TO 39, 0 TO 29) := (
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" )
);

CONSTANT B5 : ImageMatrix(0 TO 39, 0 TO 29) := (
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" )
);

--Numero 6

CONSTANT R6 : ImageMatrix(0 TO 39, 0 TO 29) := (
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" )
);

CONSTANT G6: ImageMatrix(0 TO 39, 0 TO 29) := (
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" )
);

CONSTANT B6 : ImageMatrix(0 TO 39, 0 TO 29) := (
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" )
);

--Numero 7

CONSTANT R7 : ImageMatrix(0 TO 39, 0 TO 29) := (
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" )
);

CONSTANT G7 : ImageMatrix(0 TO 39, 0 TO 29) := (
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" )
);

CONSTANT B7 : ImageMatrix(0 TO 39, 0 TO 29) := (
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" )
);

--Numero 8

CONSTANT R8 : ImageMatrix(0 TO 39, 0 TO 29) := (
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" )
);

CONSTANT G8 : ImageMatrix(0 TO 39, 0 TO 29) := (
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" )
);

CONSTANT B8 : ImageMatrix(0 TO 39, 0 TO 29) := (
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" )
);

--Numero 9 

CONSTANT R9 : ImageMatrix(0 TO 39, 0 TO 29) := (
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"00" , x"00" , x"00" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" )
);

CONSTANT G9 : ImageMatrix(0 TO 39, 0 TO 29) := (
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"00" , x"00" , x"00" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" )
);

CONSTANT B9 : ImageMatrix(0 TO 39, 0 TO 29) := (
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"00" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"00" , x"00" , x"00" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" )
);

--------------------Bars

CONSTANT BACKGROUNDBAR_R : ImageMatrix(0 TO 24, 0 TO 199) := (
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" )
);

CONSTANT BACKGROUNDBAR_G : ImageMatrix(0 TO 24, 0 TO 199) := (
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" )
);

CONSTANT BACKGROUNDBAR_B : ImageMatrix(0 TO 24, 0 TO 199) := (
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" )
);


--BoostBlue
---------------------------------------------------------------------------------------------------------------------------------------------------------------
CONSTANT CARGA_P1R : ImageMatrix(0 TO 21, 0 TO 179) := (
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" )
);

CONSTANT CARGA_P1G : ImageMatrix(0 TO 21, 0 TO 179) := (
( x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" ),
( x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" ),
( x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" ),
( x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" ),
( x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" ),
( x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" ),
( x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" ),
( x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" ),
( x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" ),
( x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" ),
( x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" ),
( x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" ),
( x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" ),
( x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" ),
( x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" ),
( x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" ),
( x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" ),
( x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" ),
( x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" ),
( x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" ),
( x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" ),
( x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" , x"A2" )
);

CONSTANT CARGA_P1B : ImageMatrix(0 TO 21, 0 TO 179) := (
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" )
);



--BoostRed
---------------------------------------------------------------------------------------------------------------------------------------------------------------

CONSTANT CARGA_P2R : ImageMatrix(0 TO 21, 0 TO 179) := (
( x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" ),
( x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" ),
( x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" ),
( x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" ),
( x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" ),
( x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" ),
( x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" ),
( x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" ),
( x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" ),
( x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" ),
( x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" ),
( x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" ),
( x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" ),
( x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" ),
( x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" ),
( x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" ),
( x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" ),
( x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" ),
( x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" ),
( x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" ),
( x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" ),
( x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" )
);

CONSTANT CARGA_P2G : ImageMatrix(0 TO 21, 0 TO 179) := (
( x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" ),
( x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" ),
( x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" ),
( x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" ),
( x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" ),
( x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" ),
( x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" ),
( x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" ),
( x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" ),
( x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" ),
( x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" ),
( x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" ),
( x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" ),
( x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" ),
( x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" ),
( x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" ),
( x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" ),
( x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" ),
( x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" ),
( x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" ),
( x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" ),
( x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" )
);

CONSTANT CARGA_P2B : ImageMatrix(0 TO 21, 0 TO 179) := (
( x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" ),
( x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" ),
( x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" ),
( x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" ),
( x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" ),
( x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" ),
( x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" ),
( x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" ),
( x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" ),
( x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" ),
( x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" ),
( x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" ),
( x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" ),
( x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" ),
( x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" ),
( x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" ),
( x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" ),
( x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" ),
( x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" ),
( x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" ),
( x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" ),
( x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" )
);


---WIN MESSAGE

CONSTANT P1winsR : ImageMatrix(0 TO 99, 0 TO 199) := (
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B3" , x"A1" , x"97" , x"91" , x"8B" , x"8B" , x"8B" , x"8C" , x"92" , x"96" , x"A1" , x"B2" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"8D" , x"71" , x"6E" , x"6E" , x"6E" , x"6E" , x"6E" , x"6E" , x"6E" , x"6E" , x"6E" , x"6E" , x"6E" , x"6E" , x"6E" , x"6E" , x"6F" , x"79" , x"7F" , x"8B" , x"A2" , x"B4" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B3" , x"95" , x"73" , x"6E" , x"6E" , x"73" , x"98" , x"B5" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B6" , x"9D" , x"75" , x"6E" , x"6E" , x"6E" , x"6E" , x"92" , x"B4" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"AA" , x"7B" , x"6E" , x"6E" , x"6F" , x"8C" , x"B2" , x"B7" , x"B7" , x"B7" , x"99" , x"74" , x"6E" , x"6E" , x"6E" , x"9E" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"A7" , x"7D" , x"6E" , x"6E" , x"6E" , x"73" , x"A3" , x"B6" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"A1" , x"79" , x"6E" , x"6E" , x"72" , x"98" , x"B5" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"AD" , x"8B" , x"69" , x"43" , x"2D" , x"22" , x"17" , x"16" , x"16" , x"18" , x"24" , x"2C" , x"41" , x"69" , x"88" , x"A6" , x"B6" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"55" , x"15" , x"0B" , x"0B" , x"0B" , x"0B" , x"0B" , x"0B" , x"0B" , x"0B" , x"0B" , x"0B" , x"0B" , x"0B" , x"0B" , x"0B" , x"0E" , x"16" , x"1C" , x"27" , x"40" , x"69" , x"9C" , x"B5" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"97" , x"5B" , x"50" , x"6C" , x"A4" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B3" , x"78" , x"1D" , x"0C" , x"0B" , x"12" , x"67" , x"B1" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B5" , x"69" , x"18" , x"0B" , x"0B" , x"0B" , x"0B" , x"46" , x"A1" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B6" , x"86" , x"22" , x"0B" , x"0B" , x"13" , x"5C" , x"AC" , x"B7" , x"B7" , x"B7" , x"71" , x"1B" , x"0B" , x"0B" , x"0B" , x"7D" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"92" , x"2F" , x"0B" , x"0B" , x"0B" , x"12" , x"60" , x"AB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"85" , x"26" , x"0C" , x"0B" , x"16" , x"70" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B4" , x"94" , x"59" , x"28" , x"10" , x"06" , x"03" , x"01" , x"00" , x"00" , x"00" , x"01" , x"02" , x"03" , x"06" , x"10" , x"25" , x"4D" , x"89" , x"B1" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"4F" , x"0A" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"01" , x"01" , x"03" , x"0D" , x"2A" , x"6F" , x"AA" , x"B6" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B6" , x"A4" , x"49" , x"07" , x"02" , x"33" , x"96" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"8A" , x"25" , x"01" , x"00" , x"01" , x"43" , x"A1" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B3" , x"40" , x"06" , x"00" , x"00" , x"00" , x"00" , x"1E" , x"8A" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B3" , x"5B" , x"0C" , x"00" , x"00" , x"14" , x"74" , x"B0" , x"B7" , x"B7" , x"B7" , x"6C" , x"11" , x"00" , x"00" , x"00" , x"79" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"90" , x"26" , x"00" , x"00" , x"00" , x"01" , x"1B" , x"76" , x"AF" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"81" , x"1C" , x"01" , x"00" , x"0B" , x"6B" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"AE" , x"71" , x"2A" , x"09" , x"01" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"01" , x"06" , x"22" , x"66" , x"A7" , x"B6" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"4F" , x"0A" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"02" , x"14" , x"63" , x"A6" , x"B6" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"A6" , x"5B" , x"13" , x"01" , x"00" , x"32" , x"95" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"9D" , x"3E" , x"04" , x"00" , x"00" , x"27" , x"8F" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"A4" , x"25" , x"01" , x"00" , x"00" , x"00" , x"00" , x"09" , x"74" , x"B4" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B1" , x"3E" , x"06" , x"00" , x"01" , x"28" , x"9A" , x"B6" , x"B7" , x"B7" , x"B7" , x"6C" , x"11" , x"00" , x"00" , x"00" , x"79" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"90" , x"26" , x"00" , x"00" , x"00" , x"00" , x"04" , x"37" , x"92" , x"B5" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"81" , x"1C" , x"01" , x"00" , x"0B" , x"6B" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B3" , x"76" , x"20" , x"04" , x"00" , x"00" , x"01" , x"06" , x"12" , x"1D" , x"30" , x"34" , x"34" , x"2E" , x"1F" , x"13" , x"06" , x"00" , x"00" , x"00" , x"01" , x"16" , x"67" , x"A9" , x"B6" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"4F" , x"0A" , x"00" , x"00" , x"07" , x"32" , x"4E" , x"51" , x"51" , x"51" , x"51" , x"51" , x"51" , x"51" , x"51" , x"51" , x"4B" , x"31" , x"1D" , x"08" , x"00" , x"00" , x"00" , x"01" , x"21" , x"7B" , x"B1" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"A4" , x"64" , x"1D" , x"02" , x"00" , x"00" , x"32" , x"95" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B0" , x"5C" , x"0A" , x"00" , x"00" , x"13" , x"82" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"79" , x"12" , x"00" , x"00" , x"04" , x"01" , x"00" , x"01" , x"4C" , x"A9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"A9" , x"27" , x"01" , x"00" , x"02" , x"43" , x"A5" , x"B7" , x"B7" , x"B7" , x"B7" , x"6C" , x"11" , x"00" , x"00" , x"00" , x"79" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"90" , x"26" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"56" , x"A6" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"81" , x"1C" , x"01" , x"00" , x"0B" , x"6B" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"96" , x"34" , x"04" , x"00" , x"00" , x"01" , x"24" , x"55" , x"6E" , x"80" , x"9E" , x"A4" , x"A4" , x"9A" , x"82" , x"6F" , x"50" , x"1C" , x"03" , x"00" , x"00" , x"01" , x"25" , x"80" , x"B2" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"4F" , x"0A" , x"00" , x"00" , x"0F" , x"6C" , x"A6" , x"AE" , x"AE" , x"AE" , x"AE" , x"AE" , x"AE" , x"AE" , x"AE" , x"AE" , x"AA" , x"95" , x"85" , x"58" , x"11" , x"01" , x"00" , x"00" , x"05" , x"3E" , x"9A" , x"B6" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B6" , x"A2" , x"52" , x"16" , x"03" , x"00" , x"00" , x"00" , x"32" , x"95" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B6" , x"74" , x"15" , x"00" , x"00" , x"05" , x"6D" , x"B4" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"59" , x"07" , x"00" , x"00" , x"22" , x"0A" , x"00" , x"00" , x"29" , x"9F" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"88" , x"16" , x"00" , x"00" , x"04" , x"62" , x"AC" , x"B7" , x"B7" , x"B7" , x"B7" , x"6C" , x"11" , x"00" , x"00" , x"00" , x"79" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"90" , x"26" , x"00" , x"00" , x"00" , x"00" , x"00" , x"01" , x"18" , x"7E" , x"B4" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"81" , x"1C" , x"01" , x"00" , x"0B" , x"6B" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B1" , x"64" , x"10" , x"00" , x"00" , x"03" , x"37" , x"83" , x"AA" , x"B1" , x"B3" , x"B6" , x"B7" , x"B7" , x"B6" , x"B3" , x"B1" , x"A6" , x"7F" , x"29" , x"04" , x"00" , x"00" , x"06" , x"46" , x"9F" , x"B6" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"4F" , x"0A" , x"00" , x"00" , x"10" , x"71" , x"AF" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"AE" , x"69" , x"1B" , x"02" , x"00" , x"00" , x"14" , x"71" , x"B1" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B6" , x"AD" , x"83" , x"39" , x"09" , x"01" , x"00" , x"00" , x"00" , x"00" , x"32" , x"95" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"90" , x"28" , x"00" , x"00" , x"00" , x"43" , x"A7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"9F" , x"34" , x"01" , x"00" , x"0F" , x"5B" , x"1B" , x"01" , x"00" , x"0B" , x"8D" , x"B5" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"63" , x"0B" , x"00" , x"00" , x"13" , x"91" , x"B6" , x"B7" , x"B7" , x"B7" , x"B7" , x"6C" , x"11" , x"00" , x"00" , x"00" , x"79" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"90" , x"26" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"01" , x"2C" , x"97" , x"B5" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"81" , x"1C" , x"01" , x"00" , x"0B" , x"6B" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"95" , x"34" , x"03" , x"00" , x"01" , x"2A" , x"8C" , x"B5" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B6" , x"8A" , x"2C" , x"04" , x"00" , x"00" , x"18" , x"79" , x"B4" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"4F" , x"0A" , x"00" , x"00" , x"10" , x"71" , x"AF" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"A4" , x"54" , x"0B" , x"00" , x"00" , x"05" , x"54" , x"AA" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B6" , x"92" , x"5F" , x"25" , x"07" , x"01" , x"00" , x"00" , x"00" , x"00" , x"00" , x"32" , x"95" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B1" , x"45" , x"02" , x"00" , x"00" , x"29" , x"9F" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"85" , x"20" , x"00" , x"00" , x"24" , x"84" , x"35" , x"04" , x"00" , x"04" , x"5D" , x"AB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B3" , x"48" , x"04" , x"00" , x"00" , x"2A" , x"9F" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"6C" , x"11" , x"00" , x"00" , x"00" , x"79" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"90" , x"26" , x"00" , x"00" , x"00" , x"06" , x"02" , x"00" , x"00" , x"08" , x"54" , x"A4" , x"B6" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"81" , x"1C" , x"01" , x"00" , x"0B" , x"6B" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"85" , x"20" , x"01" , x"00" , x"09" , x"60" , x"AE" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"AD" , x"62" , x"11" , x"00" , x"00" , x"06" , x"5D" , x"AE" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"4F" , x"0A" , x"00" , x"00" , x"10" , x"71" , x"AF" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B6" , x"82" , x"1D" , x"01" , x"00" , x"01" , x"39" , x"9B" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B3" , x"98" , x"71" , x"33" , x"11" , x"03" , x"00" , x"00" , x"05" , x"06" , x"01" , x"00" , x"00" , x"32" , x"95" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"5E" , x"09" , x"00" , x"00" , x"11" , x"98" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"6F" , x"11" , x"00" , x"01" , x"45" , x"9F" , x"53" , x"0B" , x"00" , x"01" , x"3B" , x"A3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"9C" , x"2F" , x"00" , x"00" , x"00" , x"4E" , x"AA" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"6C" , x"11" , x"00" , x"00" , x"00" , x"79" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"90" , x"26" , x"00" , x"00" , x"00" , x"29" , x"13" , x"01" , x"00" , x"01" , x"1C" , x"76" , x"B1" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"81" , x"1C" , x"01" , x"00" , x"0B" , x"6B" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"7B" , x"16" , x"00" , x"00" , x"13" , x"74" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B6" , x"88" , x"27" , x"01" , x"00" , x"01" , x"41" , x"A2" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"4F" , x"0A" , x"00" , x"00" , x"10" , x"71" , x"AF" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"91" , x"2B" , x"03" , x"00" , x"00" , x"27" , x"8D" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"9C" , x"49" , x"15" , x"04" , x"01" , x"00" , x"01" , x"0C" , x"45" , x"3E" , x"06" , x"00" , x"00" , x"32" , x"95" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"81" , x"14" , x"00" , x"00" , x"04" , x"73" , x"B0" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"A7" , x"4D" , x"06" , x"00" , x"0A" , x"64" , x"AF" , x"84" , x"16" , x"00" , x"00" , x"20" , x"8C" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"7F" , x"1C" , x"00" , x"00" , x"09" , x"76" , x"B6" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"6C" , x"11" , x"00" , x"00" , x"00" , x"79" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"90" , x"26" , x"00" , x"00" , x"00" , x"43" , x"4A" , x"0E" , x"00" , x"00" , x"04" , x"33" , x"8F" , x"B5" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"81" , x"1C" , x"01" , x"00" , x"0B" , x"6B" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"79" , x"13" , x"00" , x"00" , x"11" , x"70" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"9C" , x"3F" , x"13" , x"1B" , x"1D" , x"50" , x"A4" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"4F" , x"0A" , x"00" , x"00" , x"10" , x"71" , x"AF" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"92" , x"2F" , x"03" , x"00" , x"00" , x"22" , x"89" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"92" , x"2F" , x"03" , x"00" , x"01" , x"0B" , x"2C" , x"6D" , x"A1" , x"5F" , x"08" , x"00" , x"00" , x"32" , x"95" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"AB" , x"29" , x"01" , x"00" , x"02" , x"4E" , x"A7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"90" , x"2C" , x"02" , x"00" , x"1B" , x"7B" , x"B3" , x"9C" , x"2E" , x"04" , x"00" , x"0E" , x"67" , x"AE" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B5" , x"67" , x"0E" , x"00" , x"00" , x"1E" , x"8B" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"6C" , x"11" , x"00" , x"00" , x"00" , x"79" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"90" , x"26" , x"00" , x"00" , x"00" , x"4A" , x"8D" , x"41" , x"09" , x"00" , x"00" , x"08" , x"4E" , x"A4" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"81" , x"1C" , x"01" , x"00" , x"0B" , x"6B" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"81" , x"1D" , x"01" , x"00" , x"04" , x"4B" , x"A5" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B3" , x"A1" , x"99" , x"9C" , x"9C" , x"A6" , x"B4" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"4F" , x"0A" , x"00" , x"00" , x"10" , x"71" , x"AF" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"90" , x"2A" , x"03" , x"00" , x"00" , x"2B" , x"90" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"92" , x"2F" , x"03" , x"09" , x"29" , x"59" , x"90" , x"AE" , x"B6" , x"62" , x"08" , x"00" , x"00" , x"32" , x"95" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B3" , x"41" , x"06" , x"00" , x"01" , x"36" , x"A2" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B6" , x"7B" , x"18" , x"01" , x"01" , x"33" , x"97" , x"B6" , x"A5" , x"46" , x"07" , x"00" , x"06" , x"4F" , x"AA" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"A7" , x"4B" , x"06" , x"00" , x"00" , x"3F" , x"9F" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"6C" , x"11" , x"00" , x"00" , x"00" , x"79" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"90" , x"26" , x"00" , x"00" , x"00" , x"4B" , x"A6" , x"83" , x"25" , x"01" , x"00" , x"01" , x"15" , x"72" , x"B1" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"81" , x"1C" , x"01" , x"00" , x"0B" , x"6B" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"90" , x"2E" , x"02" , x"00" , x"01" , x"17" , x"69" , x"A7" , x"B6" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"4F" , x"0A" , x"00" , x"00" , x"10" , x"71" , x"AF" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B4" , x"7E" , x"1B" , x"01" , x"00" , x"00" , x"43" , x"A1" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"92" , x"3A" , x"2F" , x"62" , x"8B" , x"A9" , x"B4" , x"B7" , x"B7" , x"62" , x"08" , x"00" , x"00" , x"32" , x"95" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B4" , x"5F" , x"0E" , x"00" , x"00" , x"20" , x"90" , x"B4" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"AC" , x"59" , x"0B" , x"00" , x"06" , x"50" , x"A9" , x"B7" , x"B1" , x"6B" , x"11" , x"01" , x"01" , x"33" , x"97" , x"B6" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"94" , x"31" , x"03" , x"00" , x"08" , x"60" , x"AF" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"6C" , x"11" , x"00" , x"00" , x"00" , x"79" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"90" , x"26" , x"00" , x"00" , x"00" , x"4B" , x"A9" , x"AA" , x"5D" , x"0F" , x"00" , x"00" , x"01" , x"2C" , x"97" , x"B5" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"81" , x"1C" , x"01" , x"00" , x"0B" , x"6B" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"AB" , x"53" , x"09" , x"00" , x"00" , x"02" , x"18" , x"4E" , x"77" , x"A1" , x"B6" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"4F" , x"0A" , x"00" , x"00" , x"10" , x"71" , x"AF" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"A2" , x"49" , x"09" , x"00" , x"00" , x"07" , x"5D" , x"AF" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"AC" , x"96" , x"9A" , x"B0" , x"B6" , x"B7" , x"B7" , x"B7" , x"B7" , x"62" , x"08" , x"00" , x"00" , x"32" , x"95" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B6" , x"8D" , x"1F" , x"01" , x"00" , x"11" , x"6F" , x"AF" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"A0" , x"38" , x"05" , x"00" , x"11" , x"6C" , x"AE" , x"B7" , x"B7" , x"87" , x"22" , x"01" , x"00" , x"17" , x"76" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"85" , x"20" , x"01" , x"00" , x"17" , x"76" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"6C" , x"11" , x"00" , x"00" , x"00" , x"79" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"90" , x"26" , x"00" , x"00" , x"00" , x"4B" , x"A9" , x"B6" , x"A5" , x"42" , x"04" , x"00" , x"00" , x"06" , x"4F" , x"A4" , x"B6" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"81" , x"1C" , x"01" , x"00" , x"0B" , x"6B" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B6" , x"91" , x"2E" , x"03" , x"00" , x"00" , x"01" , x"06" , x"14" , x"2B" , x"4B" , x"6B" , x"8E" , x"A6" , x"AC" , x"B1" , x"B6" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"4F" , x"0A" , x"00" , x"00" , x"10" , x"71" , x"AF" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"A4" , x"56" , x"13" , x"01" , x"00" , x"01" , x"20" , x"80" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"62" , x"08" , x"00" , x"00" , x"32" , x"95" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"A0" , x"35" , x"04" , x"00" , x"08" , x"55" , x"AB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B6" , x"8F" , x"20" , x"01" , x"00" , x"21" , x"8E" , x"B4" , x"B7" , x"B7" , x"9C" , x"3C" , x"04" , x"00" , x"08" , x"5D" , x"AD" , x"B7" , x"B7" , x"B7" , x"B7" , x"B3" , x"70" , x"11" , x"00" , x"01" , x"2E" , x"90" , x"B5" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"6C" , x"11" , x"00" , x"00" , x"00" , x"79" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"90" , x"26" , x"00" , x"00" , x"00" , x"4B" , x"A9" , x"B7" , x"B7" , x"87" , x"20" , x"02" , x"00" , x"01" , x"16" , x"6C" , x"AC" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"81" , x"1C" , x"01" , x"00" , x"0B" , x"6B" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B3" , x"7D" , x"29" , x"06" , x"00" , x"00" , x"00" , x"00" , x"01" , x"06" , x"0F" , x"1B" , x"2E" , x"44" , x"67" , x"88" , x"98" , x"A7" , x"B5" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"4F" , x"0A" , x"00" , x"00" , x"10" , x"71" , x"AF" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B6" , x"9C" , x"8B" , x"79" , x"4B" , x"11" , x"01" , x"00" , x"00" , x"07" , x"4E" , x"A4" , x"B6" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"62" , x"08" , x"00" , x"00" , x"32" , x"95" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"A9" , x"4F" , x"09" , x"00" , x"02" , x"3F" , x"A3" , x"B6" , x"B7" , x"B7" , x"B7" , x"B5" , x"67" , x"10" , x"00" , x"01" , x"3E" , x"A2" , x"B7" , x"B7" , x"B7" , x"AF" , x"59" , x"09" , x"00" , x"01" , x"3B" , x"9C" , x"B7" , x"B7" , x"B7" , x"B7" , x"A6" , x"4C" , x"09" , x"00" , x"05" , x"4A" , x"A6" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"6C" , x"11" , x"00" , x"00" , x"00" , x"79" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"90" , x"26" , x"00" , x"00" , x"00" , x"4B" , x"A9" , x"B7" , x"B7" , x"AE" , x"63" , x"13" , x"01" , x"00" , x"03" , x"2F" , x"8C" , x"B5" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"81" , x"1C" , x"01" , x"00" , x"0B" , x"6B" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"AE" , x"7E" , x"3B" , x"0E" , x"01" , x"00" , x"00" , x"00" , x"00" , x"00" , x"01" , x"04" , x"07" , x"0F" , x"1C" , x"32" , x"4E" , x"74" , x"94" , x"AF" , x"B6" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"4F" , x"0A" , x"00" , x"00" , x"07" , x"31" , x"4B" , x"4F" , x"4F" , x"4F" , x"4F" , x"4F" , x"4F" , x"4F" , x"4F" , x"4F" , x"36" , x"27" , x"17" , x"09" , x"01" , x"00" , x"00" , x"01" , x"28" , x"89" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"62" , x"08" , x"00" , x"00" , x"32" , x"95" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B3" , x"72" , x"14" , x"01" , x"00" , x"28" , x"8D" , x"B5" , x"B7" , x"B7" , x"B7" , x"B3" , x"43" , x"07" , x"00" , x"04" , x"5F" , x"AC" , x"B7" , x"B7" , x"B7" , x"B6" , x"74" , x"16" , x"00" , x"00" , x"1D" , x"8B" , x"B7" , x"B7" , x"B7" , x"B7" , x"9D" , x"32" , x"04" , x"00" , x"0D" , x"61" , x"AD" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"6C" , x"11" , x"00" , x"00" , x"00" , x"79" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"90" , x"26" , x"00" , x"00" , x"00" , x"4B" , x"A9" , x"B7" , x"B7" , x"B7" , x"9D" , x"3E" , x"06" , x"00" , x"00" , x"09" , x"4D" , x"A3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"81" , x"1C" , x"01" , x"00" , x"0B" , x"6B" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B1" , x"96" , x"66" , x"2B" , x"08" , x"01" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"01" , x"04" , x"08" , x"16" , x"31" , x"5D" , x"97" , x"B4" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"4F" , x"0A" , x"00" , x"00" , x"00" , x"01" , x"01" , x"01" , x"01" , x"01" , x"01" , x"01" , x"01" , x"01" , x"01" , x"01" , x"01" , x"01" , x"00" , x"00" , x"00" , x"00" , x"04" , x"27" , x"8B" , x"B2" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"62" , x"08" , x"00" , x"00" , x"32" , x"95" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"8D" , x"27" , x"02" , x"00" , x"14" , x"73" , x"B2" , x"B7" , x"B7" , x"B7" , x"9F" , x"22" , x"01" , x"00" , x"0D" , x"8D" , x"B5" , x"B7" , x"B7" , x"B7" , x"B7" , x"92" , x"29" , x"00" , x"00" , x"07" , x"75" , x"B5" , x"B7" , x"B7" , x"B6" , x"90" , x"1C" , x"01" , x"00" , x"1D" , x"8A" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"6C" , x"11" , x"00" , x"00" , x"00" , x"79" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"90" , x"26" , x"00" , x"00" , x"00" , x"4B" , x"A9" , x"B7" , x"B7" , x"B7" , x"B3" , x"85" , x"2B" , x"03" , x"00" , x"00" , x"0E" , x"6C" , x"B1" , x"B7" , x"B7" , x"B7" , x"B7" , x"81" , x"1C" , x"01" , x"00" , x"0B" , x"6B" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B6" , x"B1" , x"9E" , x"85" , x"52" , x"2D" , x"15" , x"0A" , x"04" , x"01" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"01" , x"09" , x"28" , x"6F" , x"A6" , x"B6" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"4F" , x"0A" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"04" , x"16" , x"3C" , x"85" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"62" , x"08" , x"00" , x"00" , x"32" , x"95" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"9E" , x"3E" , x"04" , x"00" , x"09" , x"64" , x"B1" , x"B7" , x"B7" , x"B7" , x"78" , x"11" , x"00" , x"00" , x"26" , x"9F" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B1" , x"46" , x"03" , x"00" , x"01" , x"48" , x"A9" , x"B7" , x"B7" , x"B4" , x"64" , x"0E" , x"00" , x"01" , x"35" , x"A0" , x"B6" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"6C" , x"11" , x"00" , x"00" , x"00" , x"79" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"90" , x"26" , x"00" , x"00" , x"00" , x"4B" , x"A9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B1" , x"6C" , x"13" , x"00" , x"00" , x"01" , x"26" , x"8E" , x"B3" , x"B7" , x"B7" , x"B7" , x"81" , x"1C" , x"01" , x"00" , x"0B" , x"6B" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B4" , x"A9" , x"A0" , x"81" , x"5F" , x"48" , x"30" , x"1A" , x"0B" , x"03" , x"00" , x"00" , x"00" , x"00" , x"00" , x"03" , x"1A" , x"61" , x"A4" , x"B6" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"4F" , x"0A" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"07" , x"10" , x"1B" , x"2E" , x"54" , x"74" , x"99" , x"B1" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"62" , x"08" , x"00" , x"00" , x"32" , x"95" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B0" , x"5D" , x"0B" , x"00" , x"01" , x"48" , x"A4" , x"B7" , x"B7" , x"B7" , x"59" , x"07" , x"00" , x"00" , x"4B" , x"A9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"63" , x"0B" , x"00" , x"00" , x"26" , x"9E" , x"B7" , x"B7" , x"B2" , x"44" , x"07" , x"00" , x"03" , x"52" , x"A8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"6C" , x"11" , x"00" , x"00" , x"00" , x"79" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"90" , x"26" , x"00" , x"00" , x"00" , x"4B" , x"A9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"A1" , x"41" , x"05" , x"00" , x"00" , x"06" , x"4B" , x"A1" , x"B6" , x"B7" , x"B7" , x"81" , x"1C" , x"01" , x"00" , x"0B" , x"6B" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B2" , x"AC" , x"A8" , x"96" , x"7A" , x"64" , x"4D" , x"2A" , x"0D" , x"01" , x"00" , x"00" , x"00" , x"01" , x"1B" , x"74" , x"B1" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"4F" , x"0A" , x"00" , x"00" , x"0A" , x"46" , x"6C" , x"71" , x"71" , x"71" , x"71" , x"71" , x"71" , x"71" , x"71" , x"71" , x"76" , x"7D" , x"85" , x"93" , x"AB" , x"B2" , x"B6" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"62" , x"08" , x"00" , x"00" , x"32" , x"95" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B6" , x"78" , x"18" , x"00" , x"00" , x"28" , x"90" , x"B7" , x"B7" , x"A8" , x"3C" , x"01" , x"00" , x"07" , x"72" , x"B4" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"86" , x"16" , x"00" , x"00" , x"0D" , x"8B" , x"B4" , x"B7" , x"AF" , x"2A" , x"02" , x"00" , x"09" , x"82" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"6C" , x"11" , x"00" , x"00" , x"00" , x"79" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"90" , x"26" , x"00" , x"00" , x"00" , x"4B" , x"A9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B6" , x"90" , x"22" , x"02" , x"00" , x"00" , x"16" , x"6C" , x"AE" , x"B7" , x"B7" , x"81" , x"1C" , x"01" , x"00" , x"0B" , x"6B" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B6" , x"B3" , x"B1" , x"A7" , x"90" , x"77" , x"38" , x"0E" , x"01" , x"00" , x"00" , x"03" , x"32" , x"98" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"4F" , x"0A" , x"00" , x"00" , x"10" , x"71" , x"AF" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"62" , x"08" , x"00" , x"00" , x"32" , x"95" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"95" , x"2B" , x"00" , x"00" , x"13" , x"82" , x"B7" , x"B7" , x"85" , x"21" , x"00" , x"00" , x"1D" , x"89" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"AC" , x"2D" , x"03" , x"00" , x"04" , x"61" , x"AC" , x"B7" , x"85" , x"15" , x"00" , x"00" , x"20" , x"9C" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"6C" , x"11" , x"00" , x"00" , x"00" , x"79" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"90" , x"26" , x"00" , x"00" , x"00" , x"4B" , x"A9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B3" , x"69" , x"14" , x"01" , x"00" , x"01" , x"26" , x"82" , x"B3" , x"B7" , x"81" , x"1C" , x"01" , x"00" , x"0B" , x"6B" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B6" , x"A1" , x"6C" , x"22" , x"03" , x"00" , x"00" , x"07" , x"6E" , x"B1" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"4F" , x"0A" , x"00" , x"00" , x"10" , x"71" , x"AF" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"62" , x"08" , x"00" , x"00" , x"32" , x"95" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B2" , x"47" , x"03" , x"00" , x"04" , x"6B" , x"B3" , x"B7" , x"6E" , x"11" , x"00" , x"01" , x"3D" , x"9E" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B3" , x"4A" , x"09" , x"00" , x"02" , x"46" , x"A6" , x"B7" , x"69" , x"0C" , x"00" , x"00" , x"3E" , x"A6" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"6C" , x"11" , x"00" , x"00" , x"00" , x"79" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"90" , x"26" , x"00" , x"00" , x"00" , x"4B" , x"A9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B6" , x"A0" , x"4B" , x"0B" , x"00" , x"00" , x"06" , x"44" , x"9F" , x"B7" , x"81" , x"1C" , x"01" , x"00" , x"0B" , x"6B" , x"B3" , x"B7" , x"B7" , x"B7" , x"B6" , x"9D" , x"8A" , x"85" , x"80" , x"8B" , x"B0" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B6" , x"A9" , x"61" , x"11" , x"00" , x"00" , x"01" , x"47" , x"A7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"4F" , x"0A" , x"00" , x"00" , x"10" , x"71" , x"AF" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"62" , x"08" , x"00" , x"00" , x"32" , x"95" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"63" , x"0A" , x"00" , x"00" , x"47" , x"A9" , x"AA" , x"50" , x"07" , x"00" , x"08" , x"5F" , x"AF" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B5" , x"6E" , x"11" , x"00" , x"01" , x"2E" , x"A1" , x"B7" , x"50" , x"05" , x"00" , x"04" , x"67" , x"B2" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"6C" , x"11" , x"00" , x"00" , x"00" , x"79" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"90" , x"26" , x"00" , x"00" , x"00" , x"4B" , x"A9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B5" , x"89" , x"2A" , x"02" , x"00" , x"00" , x"10" , x"69" , x"AF" , x"81" , x"1C" , x"01" , x"00" , x"0B" , x"6B" , x"B3" , x"B7" , x"B7" , x"B7" , x"B1" , x"60" , x"28" , x"1D" , x"18" , x"36" , x"9B" , x"B6" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B6" , x"9C" , x"2A" , x"00" , x"00" , x"00" , x"35" , x"A2" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"4F" , x"0A" , x"00" , x"00" , x"10" , x"71" , x"AF" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"62" , x"08" , x"00" , x"00" , x"32" , x"95" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"83" , x"14" , x"00" , x"00" , x"2A" , x"A0" , x"95" , x"32" , x"03" , x"00" , x"16" , x"74" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"93" , x"24" , x"02" , x"00" , x"19" , x"81" , x"9C" , x"33" , x"01" , x"00" , x"13" , x"83" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"6C" , x"11" , x"00" , x"00" , x"00" , x"79" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"90" , x"26" , x"00" , x"00" , x"00" , x"4B" , x"A9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"AE" , x"6A" , x"15" , x"00" , x"00" , x"01" , x"21" , x"8D" , x"7E" , x"1C" , x"01" , x"00" , x"0B" , x"6B" , x"B3" , x"B7" , x"B7" , x"B7" , x"B1" , x"52" , x"0B" , x"01" , x"01" , x"18" , x"7B" , x"B1" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B6" , x"41" , x"02" , x"00" , x"00" , x"2B" , x"9F" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"4F" , x"0A" , x"00" , x"00" , x"10" , x"71" , x"AF" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"62" , x"08" , x"00" , x"00" , x"32" , x"95" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"AB" , x"2A" , x"02" , x"00" , x"13" , x"95" , x"83" , x"1D" , x"01" , x"01" , x"2E" , x"92" , x"B6" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"A3" , x"41" , x"06" , x"00" , x"0E" , x"64" , x"79" , x"1E" , x"00" , x"00" , x"31" , x"96" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"6C" , x"11" , x"00" , x"00" , x"00" , x"79" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"90" , x"26" , x"00" , x"00" , x"00" , x"4B" , x"A9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"AC" , x"4E" , x"07" , x"00" , x"00" , x"04" , x"41" , x"66" , x"1B" , x"01" , x"00" , x"0B" , x"6B" , x"B3" , x"B7" , x"B7" , x"B7" , x"B3" , x"6E" , x"11" , x"00" , x"00" , x"0A" , x"56" , x"A7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B1" , x"3D" , x"02" , x"00" , x"00" , x"34" , x"A2" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"4F" , x"0A" , x"00" , x"00" , x"10" , x"71" , x"AF" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"62" , x"08" , x"00" , x"00" , x"32" , x"95" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B3" , x"46" , x"08" , x"00" , x"06" , x"74" , x"66" , x"0F" , x"00" , x"06" , x"4B" , x"A6" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"AE" , x"62" , x"0E" , x"00" , x"09" , x"56" , x"63" , x"12" , x"00" , x"04" , x"51" , x"A9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"6C" , x"11" , x"00" , x"00" , x"00" , x"79" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"90" , x"26" , x"00" , x"00" , x"00" , x"4B" , x"A9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"8E" , x"27" , x"04" , x"00" , x"00" , x"12" , x"30" , x"11" , x"01" , x"00" , x"0B" , x"6B" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"90" , x"22" , x"02" , x"00" , x"01" , x"29" , x"89" , x"B5" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"93" , x"26" , x"00" , x"00" , x"00" , x"45" , x"A7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"4F" , x"0A" , x"00" , x"00" , x"10" , x"71" , x"AF" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"62" , x"08" , x"00" , x"00" , x"32" , x"95" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B5" , x"67" , x"0F" , x"00" , x"03" , x"47" , x"3B" , x"08" , x"00" , x"0D" , x"64" , x"AE" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B6" , x"80" , x"1C" , x"01" , x"03" , x"3D" , x"48" , x"09" , x"00" , x"0F" , x"6C" , x"B1" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"6C" , x"11" , x"00" , x"00" , x"00" , x"79" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"90" , x"26" , x"00" , x"00" , x"00" , x"4B" , x"A9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B1" , x"6F" , x"17" , x"01" , x"00" , x"02" , x"09" , x"06" , x"00" , x"00" , x"0B" , x"6B" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"A4" , x"46" , x"07" , x"00" , x"00" , x"09" , x"43" , x"9E" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"AA" , x"5E" , x"0F" , x"00" , x"00" , x"06" , x"6F" , x"B1" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"4F" , x"0A" , x"00" , x"00" , x"10" , x"71" , x"AF" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"62" , x"08" , x"00" , x"00" , x"32" , x"95" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B6" , x"90" , x"20" , x"01" , x"01" , x"27" , x"1B" , x"04" , x"00" , x"1C" , x"88" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"94" , x"32" , x"03" , x"00" , x"1C" , x"22" , x"03" , x"00" , x"23" , x"85" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"6C" , x"11" , x"00" , x"00" , x"00" , x"79" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"90" , x"26" , x"00" , x"00" , x"00" , x"4B" , x"A9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"A4" , x"4D" , x"0B" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0B" , x"6B" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B3" , x"7E" , x"21" , x"02" , x"00" , x"00" , x"09" , x"3C" , x"8B" , x"AB" , x"B5" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B4" , x"A1" , x"62" , x"1B" , x"02" , x"00" , x"01" , x"2A" , x"95" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"4F" , x"0A" , x"00" , x"00" , x"10" , x"71" , x"AF" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"62" , x"08" , x"00" , x"00" , x"32" , x"95" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"A0" , x"37" , x"05" , x"01" , x"0E" , x"06" , x"01" , x"01" , x"39" , x"A1" , x"B6" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"A8" , x"4E" , x"07" , x"00" , x"0A" , x"0C" , x"01" , x"03" , x"42" , x"A3" , x"B6" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"6C" , x"11" , x"00" , x"00" , x"00" , x"79" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"90" , x"26" , x"00" , x"00" , x"00" , x"4B" , x"A9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B5" , x"8F" , x"34" , x"04" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0B" , x"6B" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"A9" , x"5D" , x"0F" , x"00" , x"00" , x"00" , x"06" , x"22" , x"51" , x"80" , x"97" , x"A4" , x"B1" , x"B6" , x"B6" , x"AE" , x"A1" , x"97" , x"7B" , x"41" , x"13" , x"02" , x"00" , x"01" , x"15" , x"6D" , x"AF" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"4F" , x"0A" , x"00" , x"00" , x"10" , x"71" , x"AF" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"62" , x"08" , x"00" , x"00" , x"32" , x"95" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"AB" , x"57" , x"0B" , x"00" , x"01" , x"00" , x"00" , x"03" , x"58" , x"AA" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B5" , x"6C" , x"11" , x"00" , x"01" , x"01" , x"00" , x"0A" , x"59" , x"AC" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"6C" , x"11" , x"00" , x"00" , x"00" , x"79" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"90" , x"26" , x"00" , x"00" , x"00" , x"4B" , x"A9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B2" , x"74" , x"18" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0B" , x"6B" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B6" , x"9C" , x"41" , x"09" , x"01" , x"00" , x"00" , x"02" , x"0A" , x"1C" , x"32" , x"48" , x"5E" , x"69" , x"69" , x"5A" , x"43" , x"2F" , x"18" , x"07" , x"01" , x"00" , x"01" , x"0E" , x"50" , x"9D" , x"B6" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"4F" , x"0A" , x"00" , x"00" , x"10" , x"71" , x"AF" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"62" , x"08" , x"00" , x"00" , x"32" , x"95" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B4" , x"77" , x"16" , x"01" , x"00" , x"00" , x"00" , x"07" , x"83" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"86" , x"21" , x"00" , x"00" , x"00" , x"00" , x"14" , x"76" , x"B1" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"6C" , x"11" , x"00" , x"00" , x"00" , x"79" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"90" , x"26" , x"00" , x"00" , x"00" , x"4B" , x"A9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"A7" , x"49" , x"06" , x"00" , x"00" , x"00" , x"00" , x"0B" , x"6B" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B5" , x"92" , x"46" , x"0E" , x"01" , x"00" , x"00" , x"00" , x"01" , x"04" , x"06" , x"09" , x"0A" , x"0A" , x"09" , x"06" , x"04" , x"01" , x"00" , x"00" , x"00" , x"0B" , x"4E" , x"97" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"4F" , x"0A" , x"00" , x"00" , x"10" , x"71" , x"AF" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"62" , x"08" , x"00" , x"00" , x"32" , x"95" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"8D" , x"29" , x"02" , x"00" , x"00" , x"00" , x"22" , x"9C" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"AF" , x"3E" , x"01" , x"00" , x"00" , x"01" , x"2B" , x"9A" , x"B6" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"6C" , x"11" , x"00" , x"00" , x"00" , x"79" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"90" , x"26" , x"00" , x"00" , x"00" , x"4B" , x"A9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"9F" , x"31" , x"04" , x"00" , x"00" , x"00" , x"0B" , x"6B" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B6" , x"A3" , x"6F" , x"2F" , x"0E" , x"03" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"03" , x"0B" , x"2A" , x"6F" , x"A5" , x"B5" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"4F" , x"0A" , x"00" , x"00" , x"10" , x"71" , x"AF" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"62" , x"08" , x"00" , x"00" , x"32" , x"95" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"A3" , x"45" , x"05" , x"00" , x"00" , x"00" , x"43" , x"A7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"5B" , x"09" , x"00" , x"00" , x"02" , x"46" , x"A6" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"6C" , x"11" , x"00" , x"00" , x"00" , x"79" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"90" , x"26" , x"00" , x"00" , x"00" , x"4B" , x"A9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B3" , x"71" , x"1B" , x"01" , x"00" , x"00" , x"0B" , x"6B" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B6" , x"AE" , x"93" , x"67" , x"3F" , x"24" , x"16" , x"0C" , x"06" , x"01" , x"00" , x"00" , x"01" , x"07" , x"0F" , x"1E" , x"3D" , x"64" , x"90" , x"AE" , x"B6" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"80" , x"5A" , x"55" , x"55" , x"5D" , x"92" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"89" , x"59" , x"55" , x"55" , x"6F" , x"A5" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B5" , x"85" , x"59" , x"55" , x"55" , x"55" , x"87" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"8E" , x"5C" , x"55" , x"55" , x"57" , x"84" , x"B0" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"8F" , x"5E" , x"55" , x"55" , x"55" , x"96" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"A2" , x"69" , x"55" , x"55" , x"55" , x"7D" , x"AF" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"A4" , x"6F" , x"57" , x"55" , x"55" , x"5B" , x"8F" , x"B4" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B5" , x"AE" , x"A1" , x"88" , x"75" , x"67" , x"5E" , x"56" , x"55" , x"55" , x"58" , x"5F" , x"6A" , x"80" , x"A1" , x"AD" , x"B4" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B3" , x"B0" , x"AF" , x"AF" , x"B0" , x"B4" , x"B6" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B3" , x"B0" , x"AF" , x"AF" , x"B1" , x"B6" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B3" , x"B0" , x"AF" , x"AF" , x"AF" , x"B3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B4" , x"B0" , x"AF" , x"AF" , x"AF" , x"B3" , x"B6" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B4" , x"B0" , x"AF" , x"AF" , x"AF" , x"B4" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B6" , x"B1" , x"AF" , x"AF" , x"AF" , x"B3" , x"B6" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B6" , x"B2" , x"B0" , x"AF" , x"AF" , x"B0" , x"B4" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B6" , x"B4" , x"B3" , x"B1" , x"B0" , x"AF" , x"AF" , x"AF" , x"B0" , x"B1" , x"B1" , x"B3" , x"B6" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" )
);

CONSTANT P1winsG : ImageMatrix(0 TO 99, 0 TO 199) := (
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"DE" , x"D9" , x"D6" , x"D4" , x"D3" , x"D3" , x"D3" , x"D7" , x"D8" , x"DE" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"C8" , x"C5" , x"C5" , x"C5" , x"C5" , x"C5" , x"C5" , x"C5" , x"C5" , x"C5" , x"C5" , x"C5" , x"C5" , x"C5" , x"C5" , x"C6" , x"CB" , x"CD" , x"D4" , x"DF" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"D8" , x"C9" , x"C5" , x"C5" , x"C8" , x"DA" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DC" , x"C8" , x"C5" , x"C5" , x"C5" , x"C5" , x"D7" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E2" , x"CC" , x"C5" , x"C5" , x"C6" , x"D4" , x"E6" , x"E8" , x"E8" , x"E8" , x"DA" , x"C9" , x"C5" , x"C5" , x"C5" , x"DC" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E0" , x"CD" , x"C5" , x"C5" , x"C5" , x"C9" , x"DF" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DE" , x"CB" , x"C5" , x"C5" , x"C8" , x"DA" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E3" , x"D4" , x"C4" , x"B3" , x"A7" , x"A2" , x"9C" , x"9C" , x"9C" , x"9D" , x"A3" , x"A6" , x"B1" , x"C4" , x"D2" , x"E0" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"BA" , x"9B" , x"98" , x"98" , x"98" , x"98" , x"98" , x"98" , x"98" , x"98" , x"98" , x"98" , x"98" , x"98" , x"98" , x"98" , x"98" , x"9C" , x"9F" , x"A5" , x"B0" , x"C3" , x"DB" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D8" , x"BE" , x"B7" , x"C4" , x"DF" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"CB" , x"A0" , x"98" , x"98" , x"9B" , x"C2" , x"E5" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"C3" , x"9D" , x"98" , x"98" , x"98" , x"98" , x"B3" , x"DD" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D0" , x"A1" , x"97" , x"98" , x"9C" , x"BD" , x"E3" , x"E8" , x"E8" , x"E8" , x"C7" , x"A0" , x"98" , x"98" , x"98" , x"CC" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D7" , x"A9" , x"98" , x"98" , x"98" , x"9B" , x"BF" , x"E2" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D0" , x"A4" , x"97" , x"98" , x"9C" , x"C7" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"D7" , x"BC" , x"A5" , x"9A" , x"95" , x"93" , x"93" , x"92" , x"92" , x"92" , x"93" , x"93" , x"93" , x"94" , x"9A" , x"A3" , x"B5" , x"D2" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"B7" , x"97" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"93" , x"92" , x"94" , x"97" , x"A6" , x"C7" , x"E2" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"DF" , x"B4" , x"95" , x"93" , x"AB" , x"D9" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D3" , x"A3" , x"93" , x"92" , x"93" , x"B2" , x"DE" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"B0" , x"94" , x"92" , x"92" , x"92" , x"92" , x"A0" , x"D2" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"BD" , x"97" , x"92" , x"92" , x"9B" , x"C8" , x"E4" , x"E8" , x"E8" , x"E8" , x"C4" , x"9A" , x"92" , x"92" , x"92" , x"CB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"A4" , x"92" , x"92" , x"92" , x"93" , x"9F" , x"CA" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CF" , x"9F" , x"92" , x"92" , x"98" , x"C5" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E4" , x"C8" , x"A5" , x"97" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"95" , x"A2" , x"C2" , x"E1" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"B7" , x"97" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"93" , x"9B" , x"C2" , x"E0" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E0" , x"BD" , x"9B" , x"93" , x"92" , x"AA" , x"D8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DB" , x"AF" , x"93" , x"92" , x"92" , x"A4" , x"D5" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DE" , x"A3" , x"93" , x"92" , x"92" , x"92" , x"92" , x"96" , x"C8" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E5" , x"AE" , x"94" , x"92" , x"93" , x"A5" , x"DA" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"9A" , x"92" , x"92" , x"92" , x"CB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"A4" , x"92" , x"92" , x"92" , x"92" , x"94" , x"AB" , x"D8" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CF" , x"9F" , x"92" , x"92" , x"98" , x"C5" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"C9" , x"A1" , x"95" , x"92" , x"92" , x"93" , x"95" , x"9B" , x"9F" , x"A9" , x"AA" , x"AA" , x"A7" , x"A1" , x"9B" , x"95" , x"92" , x"92" , x"92" , x"92" , x"9D" , x"C2" , x"E2" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"B7" , x"97" , x"92" , x"92" , x"95" , x"AA" , x"B6" , x"B8" , x"B8" , x"B8" , x"B8" , x"B8" , x"B8" , x"B8" , x"B8" , x"B8" , x"B6" , x"AA" , x"9F" , x"95" , x"92" , x"92" , x"92" , x"93" , x"A1" , x"CD" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DE" , x"C1" , x"9F" , x"93" , x"92" , x"92" , x"AA" , x"D8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E5" , x"BD" , x"96" , x"92" , x"92" , x"9C" , x"CF" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CB" , x"9A" , x"92" , x"92" , x"93" , x"93" , x"92" , x"93" , x"B6" , x"E1" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E2" , x"A5" , x"92" , x"92" , x"93" , x"B2" , x"DF" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"9A" , x"92" , x"92" , x"92" , x"CB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"A4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"97" , x"BA" , x"E0" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CF" , x"9F" , x"92" , x"92" , x"98" , x"C5" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D9" , x"AB" , x"94" , x"92" , x"92" , x"93" , x"A3" , x"BA" , x"C5" , x"CE" , x"DC" , x"DF" , x"DF" , x"DA" , x"CF" , x"C5" , x"B8" , x"9F" , x"94" , x"92" , x"92" , x"93" , x"A3" , x"CF" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"B7" , x"97" , x"92" , x"92" , x"99" , x"C4" , x"E0" , x"E3" , x"E3" , x"E3" , x"E3" , x"E3" , x"E3" , x"E3" , x"E3" , x"E3" , x"E3" , x"D9" , x"D0" , x"BB" , x"9A" , x"92" , x"92" , x"92" , x"94" , x"AF" , x"DB" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"DE" , x"B8" , x"9C" , x"93" , x"92" , x"92" , x"92" , x"AA" , x"D8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"C8" , x"9A" , x"92" , x"92" , x"93" , x"C4" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"BC" , x"95" , x"92" , x"92" , x"A2" , x"96" , x"92" , x"92" , x"A5" , x"DD" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D2" , x"9C" , x"92" , x"92" , x"93" , x"C0" , x"E3" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"9A" , x"92" , x"92" , x"92" , x"CB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"A4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"9E" , x"CD" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CF" , x"9F" , x"92" , x"92" , x"98" , x"C5" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E5" , x"C0" , x"9A" , x"92" , x"92" , x"93" , x"AC" , x"CF" , x"E2" , x"E6" , x"E6" , x"E8" , x"E8" , x"E8" , x"E7" , x"E6" , x"E6" , x"E0" , x"CD" , x"A6" , x"93" , x"92" , x"92" , x"94" , x"B3" , x"DC" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"B7" , x"97" , x"92" , x"92" , x"99" , x"C8" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E4" , x"C4" , x"9F" , x"94" , x"92" , x"92" , x"9B" , x"C7" , x"E5" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E3" , x"CF" , x"AD" , x"97" , x"92" , x"92" , x"92" , x"92" , x"92" , x"AA" , x"D8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"A5" , x"92" , x"92" , x"92" , x"B2" , x"E0" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DC" , x"AA" , x"93" , x"92" , x"98" , x"BE" , x"9F" , x"93" , x"92" , x"98" , x"D4" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C1" , x"97" , x"92" , x"92" , x"9C" , x"D6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"9A" , x"92" , x"92" , x"92" , x"CB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"A4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A6" , x"D9" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CF" , x"9F" , x"92" , x"92" , x"98" , x"C5" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D8" , x"AB" , x"94" , x"92" , x"92" , x"A6" , x"D3" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D3" , x"A7" , x"94" , x"92" , x"92" , x"9D" , x"CB" , x"E6" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"B7" , x"97" , x"92" , x"92" , x"99" , x"C8" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DF" , x"B9" , x"98" , x"92" , x"92" , x"94" , x"B9" , x"E2" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"D7" , x"BF" , x"A3" , x"95" , x"93" , x"92" , x"92" , x"92" , x"92" , x"92" , x"AA" , x"D8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"B2" , x"93" , x"92" , x"92" , x"A6" , x"DD" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D0" , x"A1" , x"92" , x"92" , x"A2" , x"D0" , x"AB" , x"93" , x"92" , x"94" , x"BD" , x"E3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"B4" , x"94" , x"92" , x"92" , x"A6" , x"DD" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"9A" , x"92" , x"92" , x"92" , x"CB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"A4" , x"92" , x"92" , x"92" , x"95" , x"93" , x"92" , x"92" , x"96" , x"B9" , x"DF" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CF" , x"9F" , x"92" , x"92" , x"98" , x"C5" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D0" , x"A1" , x"93" , x"92" , x"96" , x"BF" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E3" , x"C1" , x"9A" , x"92" , x"92" , x"94" , x"BD" , x"E3" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"B7" , x"97" , x"92" , x"92" , x"99" , x"C8" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"CF" , x"9F" , x"92" , x"92" , x"93" , x"AD" , x"DB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"DA" , x"C7" , x"AB" , x"9A" , x"94" , x"92" , x"92" , x"94" , x"94" , x"92" , x"92" , x"92" , x"AA" , x"D8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"BE" , x"96" , x"92" , x"92" , x"9A" , x"DA" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C6" , x"9A" , x"92" , x"93" , x"B2" , x"DD" , x"BA" , x"97" , x"92" , x"93" , x"AD" , x"DF" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DB" , x"A8" , x"92" , x"92" , x"92" , x"B7" , x"E2" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"9A" , x"92" , x"92" , x"92" , x"CB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"A4" , x"92" , x"92" , x"92" , x"A6" , x"9A" , x"93" , x"92" , x"93" , x"9F" , x"CA" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CF" , x"9F" , x"92" , x"92" , x"98" , x"C5" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CC" , x"9C" , x"92" , x"92" , x"9B" , x"C8" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D2" , x"A5" , x"92" , x"92" , x"93" , x"B1" , x"DF" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"B7" , x"97" , x"92" , x"92" , x"99" , x"C8" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D7" , x"A6" , x"94" , x"92" , x"92" , x"A4" , x"D4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DB" , x"B4" , x"9B" , x"94" , x"93" , x"92" , x"93" , x"97" , x"B2" , x"AF" , x"94" , x"92" , x"92" , x"AA" , x"D8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CF" , x"9B" , x"92" , x"92" , x"93" , x"C9" , x"E5" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E0" , x"B5" , x"95" , x"92" , x"97" , x"C1" , x"E4" , x"D0" , x"9C" , x"92" , x"92" , x"A1" , x"D3" , x"E5" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CE" , x"9F" , x"92" , x"92" , x"96" , x"CA" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"9A" , x"92" , x"92" , x"92" , x"CB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"A4" , x"92" , x"92" , x"92" , x"B2" , x"B5" , x"98" , x"92" , x"92" , x"94" , x"AA" , x"D5" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CF" , x"9F" , x"92" , x"92" , x"98" , x"C5" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CB" , x"9C" , x"92" , x"92" , x"9A" , x"C7" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DB" , x"AF" , x"9B" , x"9F" , x"A0" , x"B8" , x"DF" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"B7" , x"97" , x"92" , x"92" , x"99" , x"C8" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D7" , x"A8" , x"94" , x"92" , x"92" , x"A2" , x"D3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D7" , x"A8" , x"94" , x"92" , x"92" , x"98" , x"A6" , x"C5" , x"DE" , x"BE" , x"95" , x"92" , x"92" , x"AA" , x"D8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E2" , x"A5" , x"92" , x"92" , x"93" , x"B7" , x"E0" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D6" , x"A6" , x"93" , x"92" , x"9F" , x"CC" , x"E6" , x"DB" , x"A7" , x"94" , x"92" , x"99" , x"C3" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"C3" , x"99" , x"92" , x"92" , x"A0" , x"D3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"9A" , x"92" , x"92" , x"92" , x"CB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"A4" , x"92" , x"92" , x"92" , x"B5" , x"D4" , x"B1" , x"96" , x"92" , x"92" , x"96" , x"B6" , x"DF" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CF" , x"9F" , x"92" , x"92" , x"98" , x"C5" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CF" , x"9F" , x"92" , x"92" , x"93" , x"B5" , x"DF" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"DF" , x"DA" , x"DB" , x"DC" , x"E0" , x"E6" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"B7" , x"97" , x"92" , x"92" , x"99" , x"C8" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"A6" , x"94" , x"92" , x"92" , x"A6" , x"D6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D7" , x"A8" , x"94" , x"96" , x"A5" , x"BC" , x"D5" , x"E3" , x"E7" , x"C0" , x"95" , x"92" , x"92" , x"AA" , x"D8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"B1" , x"95" , x"92" , x"93" , x"AB" , x"DE" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"CB" , x"9E" , x"92" , x"92" , x"AA" , x"D9" , x"E7" , x"DF" , x"B3" , x"95" , x"92" , x"95" , x"B7" , x"E2" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E1" , x"B5" , x"95" , x"92" , x"92" , x"B0" , x"DD" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"9A" , x"92" , x"92" , x"92" , x"CB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"A4" , x"92" , x"92" , x"92" , x"B6" , x"E1" , x"D0" , x"A4" , x"93" , x"92" , x"93" , x"9B" , x"C8" , x"E5" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CF" , x"9F" , x"92" , x"92" , x"98" , x"C5" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D6" , x"A8" , x"94" , x"92" , x"93" , x"9C" , x"C3" , x"E0" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"B7" , x"97" , x"92" , x"92" , x"99" , x"C8" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"CE" , x"9F" , x"93" , x"92" , x"92" , x"B2" , x"DE" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D7" , x"AD" , x"A8" , x"C1" , x"D3" , x"E2" , x"E6" , x"E8" , x"E8" , x"C0" , x"95" , x"92" , x"92" , x"AA" , x"D8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"BE" , x"98" , x"92" , x"92" , x"A1" , x"D6" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E2" , x"BC" , x"98" , x"92" , x"94" , x"B8" , x"E2" , x"E8" , x"E5" , x"C5" , x"9B" , x"93" , x"93" , x"AA" , x"DA" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D7" , x"A9" , x"94" , x"92" , x"96" , x"BF" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"9A" , x"92" , x"92" , x"92" , x"CB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"A4" , x"92" , x"92" , x"92" , x"B6" , x"E2" , x"E3" , x"BE" , x"99" , x"92" , x"92" , x"93" , x"A6" , x"D9" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CF" , x"9F" , x"92" , x"92" , x"98" , x"C5" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E3" , x"B9" , x"95" , x"92" , x"92" , x"94" , x"9E" , x"B6" , x"CA" , x"DE" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"B7" , x"97" , x"92" , x"92" , x"99" , x"C8" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DF" , x"B5" , x"97" , x"92" , x"92" , x"95" , x"BD" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E3" , x"D8" , x"DA" , x"E5" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"C0" , x"95" , x"92" , x"92" , x"AA" , x"D8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"D4" , x"A1" , x"92" , x"92" , x"9A" , x"C5" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DD" , x"AD" , x"94" , x"92" , x"9A" , x"C4" , x"E4" , x"E8" , x"E8" , x"D1" , x"A2" , x"93" , x"92" , x"9D" , x"CA" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D1" , x"A1" , x"93" , x"92" , x"9C" , x"C9" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"9A" , x"92" , x"92" , x"92" , x"CB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"A4" , x"92" , x"92" , x"92" , x"B6" , x"E2" , x"E7" , x"DF" , x"B1" , x"93" , x"92" , x"92" , x"95" , x"B7" , x"DE" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CF" , x"9F" , x"92" , x"92" , x"98" , x"C5" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"D7" , x"A7" , x"93" , x"92" , x"92" , x"92" , x"95" , x"9A" , x"A7" , x"B5" , x"C5" , x"D4" , x"DF" , x"E2" , x"E5" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"B7" , x"97" , x"92" , x"92" , x"99" , x"C8" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DF" , x"BA" , x"9B" , x"92" , x"92" , x"92" , x"A1" , x"CF" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C0" , x"95" , x"92" , x"92" , x"AA" , x"D8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DD" , x"AA" , x"93" , x"92" , x"96" , x"BA" , x"E3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"D5" , x"A1" , x"93" , x"92" , x"A1" , x"D4" , x"E6" , x"E8" , x"E8" , x"DB" , x"AF" , x"94" , x"92" , x"95" , x"BD" , x"E2" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"C7" , x"99" , x"92" , x"92" , x"A8" , x"D6" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"9A" , x"92" , x"92" , x"92" , x"CB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"A4" , x"92" , x"92" , x"92" , x"B6" , x"E2" , x"E8" , x"E8" , x"D1" , x"A0" , x"93" , x"92" , x"93" , x"9C" , x"C4" , x"E2" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CF" , x"9F" , x"92" , x"92" , x"98" , x"C5" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"CD" , x"A5" , x"94" , x"92" , x"92" , x"92" , x"92" , x"92" , x"95" , x"99" , x"9F" , x"A8" , x"B1" , x"C3" , x"D2" , x"DA" , x"E1" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"B7" , x"97" , x"92" , x"92" , x"99" , x"C8" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"DA" , x"D3" , x"CB" , x"B6" , x"9B" , x"93" , x"92" , x"92" , x"95" , x"B7" , x"DE" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C0" , x"95" , x"92" , x"92" , x"AA" , x"D8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E2" , x"B7" , x"96" , x"92" , x"94" , x"B0" , x"DF" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"C2" , x"99" , x"92" , x"92" , x"AE" , x"DE" , x"E8" , x"E8" , x"E8" , x"E5" , x"BC" , x"96" , x"92" , x"92" , x"AE" , x"DB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E0" , x"B5" , x"96" , x"92" , x"94" , x"B5" , x"E0" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"9A" , x"92" , x"92" , x"92" , x"CB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"A4" , x"92" , x"92" , x"92" , x"B6" , x"E2" , x"E8" , x"E8" , x"E4" , x"C1" , x"9C" , x"92" , x"92" , x"94" , x"A8" , x"D4" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CF" , x"9F" , x"92" , x"92" , x"98" , x"C5" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E4" , x"CD" , x"AE" , x"99" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"93" , x"95" , x"95" , x"99" , x"9F" , x"AA" , x"B6" , x"C8" , x"D7" , x"E5" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"B7" , x"97" , x"92" , x"92" , x"96" , x"A9" , x"B6" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"AA" , x"A4" , x"9C" , x"96" , x"93" , x"92" , x"92" , x"93" , x"A5" , x"D3" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C0" , x"95" , x"92" , x"92" , x"AA" , x"D8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"C7" , x"9A" , x"92" , x"92" , x"A4" , x"D4" , x"E7" , x"E8" , x"E8" , x"E8" , x"E7" , x"B2" , x"95" , x"92" , x"94" , x"BF" , x"E2" , x"E8" , x"E8" , x"E8" , x"E7" , x"C8" , x"9C" , x"92" , x"92" , x"9F" , x"D3" , x"E8" , x"E8" , x"E8" , x"E8" , x"DC" , x"A9" , x"94" , x"92" , x"98" , x"BF" , x"E3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"9A" , x"92" , x"92" , x"92" , x"CB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"A4" , x"92" , x"92" , x"92" , x"B6" , x"E2" , x"E8" , x"E8" , x"E8" , x"DC" , x"AF" , x"95" , x"92" , x"92" , x"96" , x"B6" , x"DF" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CF" , x"9F" , x"92" , x"92" , x"98" , x"C5" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E5" , x"D8" , x"C2" , x"A7" , x"96" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"94" , x"96" , x"9C" , x"A9" , x"BD" , x"D9" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"B7" , x"97" , x"92" , x"92" , x"92" , x"92" , x"93" , x"93" , x"93" , x"93" , x"93" , x"93" , x"93" , x"93" , x"93" , x"93" , x"92" , x"93" , x"92" , x"92" , x"92" , x"92" , x"94" , x"A4" , x"D4" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C0" , x"95" , x"92" , x"92" , x"AA" , x"D8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D4" , x"A4" , x"93" , x"92" , x"9A" , x"C8" , x"E6" , x"E8" , x"E8" , x"E8" , x"DC" , x"A2" , x"93" , x"92" , x"97" , x"D4" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"D7" , x"A6" , x"92" , x"92" , x"95" , x"C9" , x"E7" , x"E8" , x"E8" , x"E7" , x"D6" , x"9F" , x"92" , x"92" , x"9F" , x"D3" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"9A" , x"92" , x"92" , x"92" , x"CB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"A4" , x"92" , x"92" , x"92" , x"B6" , x"E2" , x"E8" , x"E8" , x"E8" , x"E6" , x"D0" , x"A7" , x"94" , x"92" , x"92" , x"98" , x"C5" , x"E5" , x"E8" , x"E8" , x"E8" , x"E8" , x"CF" , x"9F" , x"92" , x"92" , x"98" , x"C5" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"E5" , x"DC" , x"D0" , x"B9" , x"A7" , x"9B" , x"97" , x"93" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"93" , x"97" , x"A5" , x"C7" , x"E0" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"B7" , x"97" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"93" , x"9C" , x"AE" , x"D1" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C0" , x"95" , x"92" , x"92" , x"AA" , x"D8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DC" , x"AF" , x"93" , x"92" , x"96" , x"C1" , x"E5" , x"E8" , x"E8" , x"E8" , x"CA" , x"9A" , x"92" , x"92" , x"A3" , x"DD" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"B3" , x"93" , x"92" , x"92" , x"B4" , x"E2" , x"E8" , x"E8" , x"E6" , x"C0" , x"98" , x"92" , x"93" , x"AB" , x"DE" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"9A" , x"92" , x"92" , x"92" , x"CB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"A4" , x"92" , x"92" , x"92" , x"B6" , x"E2" , x"E8" , x"E8" , x"E8" , x"E8" , x"E5" , x"C4" , x"9C" , x"92" , x"92" , x"92" , x"A4" , x"D5" , x"E6" , x"E8" , x"E8" , x"E8" , x"CF" , x"9F" , x"92" , x"92" , x"98" , x"C5" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"E2" , x"DD" , x"CF" , x"BE" , x"B4" , x"A9" , x"9E" , x"98" , x"94" , x"92" , x"92" , x"92" , x"92" , x"92" , x"94" , x"9D" , x"C0" , x"DE" , x"E7" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"B7" , x"97" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"96" , x"99" , x"A0" , x"A8" , x"B9" , x"C9" , x"DA" , x"E5" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C0" , x"95" , x"92" , x"92" , x"AA" , x"D8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E5" , x"BE" , x"97" , x"92" , x"93" , x"B4" , x"DF" , x"E8" , x"E8" , x"E8" , x"BC" , x"95" , x"92" , x"92" , x"B5" , x"E2" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C1" , x"97" , x"92" , x"92" , x"A4" , x"DC" , x"E8" , x"E8" , x"E6" , x"B1" , x"95" , x"92" , x"93" , x"B9" , x"E1" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"9A" , x"92" , x"92" , x"92" , x"CB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"A4" , x"92" , x"92" , x"92" , x"B6" , x"E2" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DE" , x"B1" , x"94" , x"92" , x"92" , x"94" , x"B5" , x"DD" , x"E8" , x"E8" , x"E8" , x"CF" , x"9F" , x"92" , x"92" , x"98" , x"C5" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"E2" , x"E1" , x"D8" , x"CC" , x"C1" , x"B6" , x"A7" , x"97" , x"93" , x"92" , x"92" , x"92" , x"92" , x"9F" , x"C8" , x"E5" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"B7" , x"97" , x"92" , x"92" , x"97" , x"B3" , x"C4" , x"C7" , x"C7" , x"C7" , x"C7" , x"C7" , x"C7" , x"C7" , x"C7" , x"C7" , x"C9" , x"CD" , x"D1" , x"D7" , x"E2" , x"E6" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C0" , x"95" , x"92" , x"92" , x"AA" , x"D8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"CA" , x"9E" , x"92" , x"92" , x"A5" , x"D6" , x"E8" , x"E8" , x"E1" , x"AE" , x"92" , x"92" , x"95" , x"C8" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D2" , x"9C" , x"92" , x"92" , x"98" , x"D3" , x"E6" , x"E8" , x"E4" , x"A6" , x"93" , x"92" , x"96" , x"CF" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"9A" , x"92" , x"92" , x"92" , x"CB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"A4" , x"92" , x"92" , x"92" , x"B6" , x"E2" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"D6" , x"A2" , x"93" , x"92" , x"92" , x"9D" , x"C5" , x"E4" , x"E8" , x"E8" , x"CF" , x"9F" , x"92" , x"92" , x"98" , x"C5" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"E6" , x"E5" , x"E1" , x"D6" , x"CA" , x"AC" , x"98" , x"93" , x"92" , x"92" , x"94" , x"A9" , x"D9" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"B7" , x"97" , x"92" , x"92" , x"99" , x"C8" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C0" , x"95" , x"92" , x"92" , x"AA" , x"D8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D8" , x"A7" , x"92" , x"92" , x"9B" , x"CF" , x"E8" , x"E8" , x"D1" , x"A2" , x"92" , x"92" , x"9F" , x"D3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E2" , x"A7" , x"94" , x"92" , x"94" , x"C0" , x"E2" , x"E8" , x"D0" , x"9B" , x"92" , x"92" , x"A1" , x"DB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"9A" , x"92" , x"92" , x"92" , x"CB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"A4" , x"92" , x"92" , x"92" , x"B6" , x"E2" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"C4" , x"9A" , x"92" , x"92" , x"92" , x"A4" , x"CF" , x"E7" , x"E8" , x"CF" , x"9F" , x"92" , x"92" , x"98" , x"C5" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"DE" , x"C4" , x"A2" , x"94" , x"92" , x"92" , x"95" , x"C5" , x"E6" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"B7" , x"97" , x"92" , x"92" , x"99" , x"C8" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C0" , x"95" , x"92" , x"92" , x"AA" , x"D8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"B3" , x"94" , x"92" , x"93" , x"C4" , x"E7" , x"E8" , x"C5" , x"9B" , x"92" , x"92" , x"AE" , x"DC" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"B4" , x"96" , x"92" , x"93" , x"B3" , x"DF" , x"E8" , x"C4" , x"97" , x"92" , x"92" , x"AF" , x"E0" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"9A" , x"92" , x"92" , x"92" , x"CB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"A4" , x"92" , x"92" , x"92" , x"B6" , x"E2" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DE" , x"B5" , x"98" , x"92" , x"92" , x"95" , x"B2" , x"DD" , x"E8" , x"CF" , x"9F" , x"92" , x"92" , x"98" , x"C5" , x"E7" , x"E8" , x"E8" , x"E8" , x"E7" , x"DB" , x"D3" , x"D0" , x"CF" , x"D4" , x"E5" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E1" , x"C0" , x"9A" , x"92" , x"92" , x"92" , x"B4" , x"E1" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"B7" , x"97" , x"92" , x"92" , x"99" , x"C8" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C0" , x"95" , x"92" , x"92" , x"AA" , x"D8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C1" , x"97" , x"92" , x"92" , x"B4" , x"E2" , x"E2" , x"B7" , x"96" , x"92" , x"96" , x"BF" , x"E5" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"C5" , x"9A" , x"92" , x"93" , x"A7" , x"DE" , x"E8" , x"B8" , x"94" , x"92" , x"94" , x"C2" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"9A" , x"92" , x"92" , x"92" , x"CB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"A4" , x"92" , x"92" , x"92" , x"B6" , x"E2" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"D2" , x"A6" , x"93" , x"92" , x"92" , x"9A" , x"C3" , x"E4" , x"CF" , x"9F" , x"92" , x"92" , x"98" , x"C5" , x"E7" , x"E8" , x"E8" , x"E8" , x"E5" , x"BF" , x"A5" , x"A0" , x"9E" , x"AB" , x"DB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DB" , x"A6" , x"92" , x"92" , x"92" , x"AB" , x"DF" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"B7" , x"97" , x"92" , x"92" , x"99" , x"C8" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C0" , x"95" , x"92" , x"92" , x"AA" , x"D8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CF" , x"9B" , x"92" , x"92" , x"A7" , x"DE" , x"D7" , x"AA" , x"94" , x"92" , x"9C" , x"C8" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D8" , x"A1" , x"93" , x"92" , x"9E" , x"CF" , x"DB" , x"AA" , x"93" , x"92" , x"9B" , x"CF" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"9A" , x"92" , x"92" , x"92" , x"CB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"A4" , x"92" , x"92" , x"92" , x"B6" , x"E2" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E4" , x"C4" , x"9B" , x"92" , x"92" , x"92" , x"A2" , x"D4" , x"CD" , x"9F" , x"92" , x"92" , x"98" , x"C5" , x"E7" , x"E8" , x"E8" , x"E8" , x"E5" , x"B8" , x"98" , x"93" , x"92" , x"9D" , x"CC" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"B0" , x"92" , x"92" , x"92" , x"A7" , x"DE" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"B7" , x"97" , x"92" , x"92" , x"99" , x"C8" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C0" , x"95" , x"92" , x"92" , x"AA" , x"D8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E2" , x"A6" , x"93" , x"92" , x"9C" , x"D9" , x"CF" , x"9F" , x"92" , x"92" , x"A7" , x"D6" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DF" , x"B1" , x"94" , x"92" , x"98" , x"C0" , x"CB" , x"A0" , x"92" , x"92" , x"A9" , x"D8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"9A" , x"92" , x"92" , x"92" , x"CB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"A4" , x"92" , x"92" , x"92" , x"B6" , x"E2" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E2" , x"B7" , x"95" , x"92" , x"92" , x"94" , x"B1" , x"C2" , x"9F" , x"92" , x"92" , x"98" , x"C5" , x"E7" , x"E8" , x"E8" , x"E8" , x"E6" , x"C5" , x"9A" , x"92" , x"92" , x"97" , x"BB" , x"E0" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E5" , x"AD" , x"93" , x"92" , x"92" , x"AA" , x"DF" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"B7" , x"97" , x"92" , x"92" , x"99" , x"C8" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C0" , x"95" , x"92" , x"92" , x"AA" , x"D8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"B2" , x"96" , x"92" , x"94" , x"C8" , x"C2" , x"99" , x"92" , x"94" , x"B6" , x"E0" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E3" , x"C1" , x"98" , x"92" , x"96" , x"BA" , x"C1" , x"9B" , x"92" , x"94" , x"B8" , x"E2" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"9A" , x"92" , x"92" , x"92" , x"CB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"A4" , x"92" , x"92" , x"92" , x"B6" , x"E2" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"A4" , x"94" , x"92" , x"92" , x"9B" , x"A9" , x"9A" , x"92" , x"92" , x"98" , x"C5" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"D6" , x"A1" , x"93" , x"92" , x"93" , x"A6" , x"D2" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D8" , x"A4" , x"92" , x"92" , x"92" , x"B2" , x"E1" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"B7" , x"97" , x"92" , x"92" , x"99" , x"C8" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C0" , x"95" , x"92" , x"92" , x"AA" , x"D8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"C2" , x"99" , x"92" , x"94" , x"B3" , x"AE" , x"96" , x"92" , x"97" , x"C1" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CF" , x"9E" , x"92" , x"94" , x"AE" , x"B4" , x"96" , x"92" , x"99" , x"C4" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"9A" , x"92" , x"92" , x"92" , x"CB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"A4" , x"92" , x"92" , x"92" , x"B6" , x"E2" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"C6" , x"9D" , x"92" , x"92" , x"94" , x"96" , x"95" , x"92" , x"92" , x"98" , x"C5" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"DE" , x"B2" , x"95" , x"92" , x"92" , x"97" , x"B2" , x"DC" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E2" , x"BE" , x"9A" , x"92" , x"92" , x"94" , x"C6" , x"E6" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"B7" , x"97" , x"92" , x"92" , x"99" , x"C8" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C0" , x"95" , x"92" , x"92" , x"AA" , x"D8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"D4" , x"A1" , x"92" , x"93" , x"A3" , x"9F" , x"94" , x"92" , x"9F" , x"D1" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D7" , x"AA" , x"94" , x"92" , x"9F" , x"A3" , x"94" , x"92" , x"A3" , x"D1" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"9A" , x"92" , x"92" , x"92" , x"CB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"A4" , x"92" , x"92" , x"92" , x"B6" , x"E2" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DF" , x"B5" , x"97" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"98" , x"C5" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E5" , x"CD" , x"A1" , x"94" , x"92" , x"92" , x"96" , x"AE" , x"D4" , x"E2" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"DD" , x"C0" , x"9F" , x"94" , x"92" , x"93" , x"A6" , x"D8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"B7" , x"97" , x"92" , x"92" , x"99" , x"C8" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C0" , x"95" , x"92" , x"92" , x"AA" , x"D8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DD" , x"AC" , x"94" , x"92" , x"99" , x"94" , x"92" , x"93" , x"AD" , x"DE" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E1" , x"B6" , x"95" , x"92" , x"97" , x"97" , x"92" , x"94" , x"B1" , x"DF" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"9A" , x"92" , x"92" , x"92" , x"CB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"A4" , x"92" , x"92" , x"92" , x"B6" , x"E2" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"D5" , x"AA" , x"94" , x"92" , x"92" , x"92" , x"92" , x"92" , x"98" , x"C5" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E2" , x"BD" , x"9A" , x"92" , x"92" , x"92" , x"94" , x"A2" , x"B8" , x"CE" , x"D9" , x"DE" , x"E5" , x"E7" , x"E7" , x"E3" , x"DE" , x"D9" , x"CC" , x"B0" , x"9B" , x"94" , x"92" , x"93" , x"9B" , x"C6" , x"E5" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"B7" , x"97" , x"92" , x"92" , x"99" , x"C8" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C0" , x"95" , x"92" , x"92" , x"AA" , x"D8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E2" , x"BB" , x"98" , x"92" , x"93" , x"92" , x"92" , x"93" , x"BC" , x"E2" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"C4" , x"99" , x"92" , x"93" , x"93" , x"92" , x"97" , x"BC" , x"E2" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"9A" , x"92" , x"92" , x"92" , x"CB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"A4" , x"92" , x"92" , x"92" , x"B6" , x"E2" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"C9" , x"9D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"98" , x"C5" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DB" , x"B0" , x"96" , x"92" , x"92" , x"92" , x"93" , x"97" , x"9F" , x"AA" , x"B4" , x"BE" , x"C3" , x"C3" , x"BD" , x"B2" , x"A8" , x"9D" , x"95" , x"92" , x"92" , x"93" , x"98" , x"B7" , x"DB" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"B7" , x"97" , x"92" , x"92" , x"99" , x"C8" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C0" , x"95" , x"92" , x"92" , x"AA" , x"D8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"CA" , x"9C" , x"92" , x"92" , x"92" , x"92" , x"94" , x"D0" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D1" , x"A1" , x"92" , x"92" , x"92" , x"92" , x"9B" , x"C9" , x"E5" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"9A" , x"92" , x"92" , x"92" , x"CB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"A4" , x"92" , x"92" , x"92" , x"B6" , x"E2" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E2" , x"B4" , x"95" , x"92" , x"92" , x"92" , x"92" , x"98" , x"C5" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"D6" , x"B3" , x"99" , x"92" , x"92" , x"92" , x"92" , x"93" , x"94" , x"95" , x"96" , x"97" , x"97" , x"96" , x"94" , x"94" , x"92" , x"92" , x"92" , x"92" , x"97" , x"B6" , x"D8" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"B7" , x"97" , x"92" , x"92" , x"99" , x"C8" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C0" , x"95" , x"92" , x"92" , x"AA" , x"D8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D4" , x"A5" , x"93" , x"92" , x"92" , x"92" , x"A3" , x"DB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E5" , x"AF" , x"93" , x"92" , x"92" , x"93" , x"A6" , x"DB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"9A" , x"92" , x"92" , x"92" , x"CB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"A4" , x"92" , x"92" , x"92" , x"B6" , x"E2" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DC" , x"A9" , x"93" , x"92" , x"92" , x"92" , x"98" , x"C5" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DF" , x"C7" , x"A8" , x"98" , x"93" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"94" , x"98" , x"A5" , x"C6" , x"DF" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"B7" , x"97" , x"92" , x"92" , x"99" , x"C8" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C0" , x"95" , x"92" , x"92" , x"AA" , x"D8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DF" , x"B2" , x"94" , x"92" , x"92" , x"92" , x"B3" , x"E1" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"BD" , x"97" , x"92" , x"92" , x"93" , x"B3" , x"DF" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"9A" , x"92" , x"92" , x"92" , x"CB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"A4" , x"92" , x"92" , x"92" , x"B6" , x"E2" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"C7" , x"9F" , x"93" , x"92" , x"92" , x"98" , x"C5" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E4" , x"D8" , x"C2" , x"AF" , x"A3" , x"9C" , x"97" , x"95" , x"92" , x"92" , x"92" , x"93" , x"95" , x"99" , x"A0" , x"AE" , x"C1" , x"D6" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CF" , x"BD" , x"B9" , x"B9" , x"BD" , x"D7" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D2" , x"BB" , x"B9" , x"B9" , x"C6" , x"E0" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"D0" , x"BC" , x"B9" , x"B9" , x"B9" , x"D1" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"BD" , x"B9" , x"B9" , x"BA" , x"D0" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"BE" , x"B9" , x"B9" , x"B9" , x"D8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DF" , x"C4" , x"B9" , x"B9" , x"B9" , x"CD" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DF" , x"C6" , x"BA" , x"B9" , x"B9" , x"BD" , x"D5" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"E3" , x"DE" , x"D2" , x"C9" , x"C3" , x"BD" , x"B9" , x"B9" , x"B9" , x"BB" , x"BF" , x"C4" , x"CE" , x"DE" , x"E3" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"E5" , x"E4" , x"E4" , x"E5" , x"E6" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"E5" , x"E4" , x"E4" , x"E6" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"E5" , x"E4" , x"E4" , x"E4" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"E5" , x"E4" , x"E4" , x"E4" , x"E6" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"E5" , x"E4" , x"E4" , x"E4" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"E5" , x"E4" , x"E4" , x"E4" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"E6" , x"E5" , x"E4" , x"E4" , x"E5" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"E7" , x"E6" , x"E4" , x"E4" , x"E4" , x"E4" , x"E5" , x"E5" , x"E6" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" )
);

CONSTANT P1winsB : ImageMatrix(0 TO 99, 0 TO 199) := (
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"95" , x"9E" , x"A3" , x"A7" , x"A9" , x"AB" , x"AB" , x"A9" , x"A6" , x"A4" , x"9E" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"A9" , x"B7" , x"BA" , x"BA" , x"BA" , x"BA" , x"BA" , x"BA" , x"BA" , x"BA" , x"BA" , x"BA" , x"BA" , x"BA" , x"BA" , x"BA" , x"B9" , x"B3" , x"AF" , x"AA" , x"9C" , x"94" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"94" , x"A5" , x"B8" , x"BA" , x"BA" , x"B7" , x"A3" , x"93" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A0" , x"B5" , x"BA" , x"BA" , x"BA" , x"BA" , x"A7" , x"94" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"99" , x"B3" , x"BA" , x"BA" , x"B9" , x"AA" , x"95" , x"92" , x"92" , x"92" , x"A2" , x"B7" , x"BA" , x"BA" , x"BA" , x"9F" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"9A" , x"B2" , x"BA" , x"BA" , x"BA" , x"B8" , x"9C" , x"93" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"9E" , x"B3" , x"BA" , x"BA" , x"B7" , x"A2" , x"93" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"97" , x"A9" , x"BC" , x"D1" , x"DC" , x"E3" , x"E8" , x"EA" , x"EA" , x"E7" , x"E2" , x"DC" , x"D2" , x"BC" , x"AC" , x"9B" , x"93" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"C6" , x"EA" , x"EF" , x"EF" , x"EF" , x"EF" , x"EF" , x"EF" , x"EF" , x"EF" , x"EF" , x"EF" , x"EF" , x"EF" , x"EF" , x"EF" , x"EE" , x"E9" , x"E5" , x"E0" , x"D2" , x"BB" , x"A1" , x"93" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A3" , x"C4" , x"C9" , x"BB" , x"9C" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"94" , x"B4" , x"E5" , x"EF" , x"EF" , x"EB" , x"BF" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"93" , x"BD" , x"E6" , x"EF" , x"EF" , x"EF" , x"EF" , x"CF" , x"9D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"AD" , x"E3" , x"EE" , x"EF" , x"EA" , x"C3" , x"98" , x"92" , x"92" , x"92" , x"B8" , x"E7" , x"EF" , x"EF" , x"EF" , x"B2" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A6" , x"DD" , x"EF" , x"EF" , x"EF" , x"EC" , x"C0" , x"98" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"AD" , x"E0" , x"EF" , x"EF" , x"E9" , x"B9" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"94" , x"A5" , x"C5" , x"DF" , x"ED" , x"F1" , x"F3" , x"F4" , x"F5" , x"F5" , x"F5" , x"F5" , x"F4" , x"F3" , x"F2" , x"ED" , x"E1" , x"CB" , x"AA" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"CA" , x"F0" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F3" , x"ED" , x"DE" , x"B9" , x"9A" , x"93" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"93" , x"9D" , x"CD" , x"F1" , x"F4" , x"DA" , x"A5" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"AA" , x"E1" , x"F4" , x"F5" , x"F5" , x"D0" , x"9D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"95" , x"D3" , x"F2" , x"F5" , x"F5" , x"F5" , x"F5" , x"E5" , x"AA" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"94" , x"C5" , x"EF" , x"F5" , x"F5" , x"EA" , x"B6" , x"95" , x"92" , x"92" , x"92" , x"BA" , x"EC" , x"F5" , x"F5" , x"F5" , x"B4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A8" , x"E1" , x"F5" , x"F5" , x"F5" , x"F5" , x"E6" , x"B5" , x"96" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"AF" , x"E5" , x"F5" , x"F5" , x"EF" , x"BB" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"97" , x"B7" , x"DE" , x"F0" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F2" , x"E3" , x"BD" , x"9A" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"CA" , x"F0" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F4" , x"EA" , x"C0" , x"9B" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"9C" , x"C4" , x"EB" , x"F5" , x"F5" , x"DB" , x"A4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"9F" , x"D3" , x"F2" , x"F5" , x"F5" , x"E0" , x"A7" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"9D" , x"E1" , x"F4" , x"F5" , x"F5" , x"F5" , x"F5" , x"F0" , x"B6" , x"93" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"95" , x"D4" , x"F2" , x"F5" , x"F5" , x"E0" , x"A3" , x"92" , x"92" , x"92" , x"92" , x"BA" , x"EC" , x"F5" , x"F5" , x"F5" , x"B4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A8" , x"E1" , x"F5" , x"F5" , x"F5" , x"F5" , x"F3" , x"D9" , x"A7" , x"93" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"AF" , x"E5" , x"F5" , x"F5" , x"EF" , x"BB" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"94" , x"B4" , x"E3" , x"F3" , x"F5" , x"F5" , x"F5" , x"F2" , x"EB" , x"E5" , x"DA" , x"D9" , x"D9" , x"DD" , x"E5" , x"EB" , x"F2" , x"F5" , x"F5" , x"F5" , x"F4" , x"E9" , x"BE" , x"9A" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"CA" , x"F0" , x"F5" , x"F5" , x"F2" , x"DA" , x"CB" , x"C9" , x"C9" , x"C9" , x"C9" , x"C9" , x"C9" , x"C9" , x"C9" , x"C9" , x"CB" , x"DB" , x"E5" , x"F0" , x"F5" , x"F5" , x"F5" , x"F5" , x"E2" , x"B3" , x"96" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"9C" , x"C0" , x"E6" , x"F4" , x"F5" , x"F5" , x"DB" , x"A4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"96" , x"C3" , x"F0" , x"F5" , x"F5" , x"EA" , x"AF" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"B4" , x"EB" , x"F5" , x"F5" , x"F2" , x"F4" , x"F5" , x"F5" , x"CC" , x"99" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"9B" , x"E0" , x"F4" , x"F5" , x"F4" , x"D1" , x"9C" , x"92" , x"92" , x"92" , x"92" , x"BA" , x"EC" , x"F5" , x"F5" , x"F5" , x"B4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A8" , x"E1" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"EE" , x"C6" , x"9B" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"AF" , x"E5" , x"F5" , x"F5" , x"EF" , x"BB" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A5" , x"D9" , x"F3" , x"F5" , x"F5" , x"F4" , x"E2" , x"C8" , x"BA" , x"B0" , x"A0" , x"9C" , x"9C" , x"A2" , x"AF" , x"B8" , x"CA" , x"E5" , x"F3" , x"F5" , x"F5" , x"F4" , x"E0" , x"AF" , x"95" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"CA" , x"F0" , x"F5" , x"F5" , x"ED" , x"BB" , x"9B" , x"97" , x"97" , x"97" , x"97" , x"97" , x"97" , x"97" , x"97" , x"97" , x"9A" , x"A5" , x"AC" , x"C5" , x"EC" , x"F5" , x"F5" , x"F5" , x"F2" , x"D4" , x"A1" , x"93" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"9D" , x"C9" , x"E8" , x"F3" , x"F5" , x"F5" , x"F5" , x"DB" , x"A4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"B6" , x"EA" , x"F5" , x"F5" , x"F2" , x"B9" , x"94" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"C5" , x"F1" , x"F5" , x"F5" , x"E1" , x"EF" , x"F5" , x"F5" , x"DF" , x"9F" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"AC" , x"E9" , x"F5" , x"F5" , x"F2" , x"C0" , x"98" , x"92" , x"92" , x"92" , x"92" , x"BA" , x"EC" , x"F5" , x"F5" , x"F5" , x"B4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A8" , x"E1" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"E8" , x"B2" , x"94" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"AF" , x"E5" , x"F5" , x"F5" , x"EF" , x"BB" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"95" , x"BF" , x"ED" , x"F5" , x"F5" , x"F3" , x"D8" , x"AD" , x"9A" , x"95" , x"94" , x"92" , x"92" , x"92" , x"93" , x"94" , x"95" , x"9B" , x"B0" , x"E0" , x"F3" , x"F5" , x"F5" , x"F1" , x"CF" , x"9F" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"CA" , x"F0" , x"F5" , x"F5" , x"ED" , x"B8" , x"96" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"98" , x"BB" , x"E7" , x"F4" , x"F5" , x"F5" , x"EA" , x"B8" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"98" , x"AF" , x"D6" , x"F0" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"DB" , x"A4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A7" , x"DF" , x"F5" , x"F5" , x"F5" , x"D1" , x"9A" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"9E" , x"D9" , x"F4" , x"F5" , x"EC" , x"C4" , x"E7" , x"F5" , x"F5" , x"EF" , x"A9" , x"93" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"BF" , x"F0" , x"F5" , x"F5" , x"EB" , x"A7" , x"93" , x"92" , x"92" , x"92" , x"92" , x"BA" , x"EC" , x"F5" , x"F5" , x"F5" , x"B4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A8" , x"E1" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"DD" , x"A4" , x"93" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"AF" , x"E5" , x"F5" , x"F5" , x"EF" , x"BB" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A4" , x"D9" , x"F3" , x"F5" , x"F5" , x"DE" , x"A9" , x"93" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"93" , x"AB" , x"DC" , x"F3" , x"F5" , x"F5" , x"E8" , x"B3" , x"94" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"CA" , x"F0" , x"F5" , x"F5" , x"ED" , x"B8" , x"96" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"9B" , x"C8" , x"EE" , x"F5" , x"F5" , x"F2" , x"C7" , x"9A" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A6" , x"C1" , x"E1" , x"F1" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"DB" , x"A4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"95" , x"CF" , x"F4" , x"F5" , x"F5" , x"DF" , x"9F" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"AD" , x"E4" , x"F5" , x"F5" , x"E3" , x"AE" , x"D8" , x"F2" , x"F5" , x"F3" , x"C2" , x"98" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"95" , x"CD" , x"F3" , x"F5" , x"F5" , x"DE" , x"9F" , x"92" , x"92" , x"92" , x"92" , x"92" , x"BA" , x"EC" , x"F5" , x"F5" , x"F5" , x"B4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A8" , x"E1" , x"F5" , x"F5" , x"F5" , x"F1" , x"F4" , x"F5" , x"F5" , x"F1" , x"C7" , x"9C" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"AF" , x"E5" , x"F5" , x"F5" , x"EF" , x"BB" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"AD" , x"E4" , x"F4" , x"F5" , x"F0" , x"C2" , x"97" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"98" , x"BF" , x"ED" , x"F5" , x"F5" , x"F2" , x"C2" , x"97" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"CA" , x"F0" , x"F5" , x"F5" , x"ED" , x"B8" , x"96" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"93" , x"AF" , x"E5" , x"F5" , x"F5" , x"F5" , x"D6" , x"A2" , x"92" , x"92" , x"92" , x"92" , x"92" , x"95" , x"A2" , x"B7" , x"DA" , x"EC" , x"F3" , x"F5" , x"F5" , x"F3" , x"F1" , x"F5" , x"F5" , x"F5" , x"DB" , x"A4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"C2" , x"F1" , x"F5" , x"F5" , x"EC" , x"A3" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"BA" , x"EC" , x"F5" , x"F4" , x"D0" , x"A0" , x"C8" , x"F0" , x"F5" , x"F4" , x"D4" , x"9C" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A1" , x"DB" , x"F5" , x"F5" , x"F5" , x"CA" , x"99" , x"92" , x"92" , x"92" , x"92" , x"92" , x"BA" , x"EC" , x"F5" , x"F5" , x"F5" , x"B4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A8" , x"E1" , x"F5" , x"F5" , x"F5" , x"E0" , x"EB" , x"F4" , x"F5" , x"F5" , x"E6" , x"B4" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"AF" , x"E5" , x"F5" , x"F5" , x"EF" , x"BB" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"B2" , x"E9" , x"F5" , x"F5" , x"EA" , x"B7" , x"94" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"AB" , x"E1" , x"F4" , x"F5" , x"F5" , x"D2" , x"9D" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"CA" , x"F0" , x"F5" , x"F5" , x"ED" , x"B8" , x"96" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A7" , x"DD" , x"F3" , x"F5" , x"F5" , x"E0" , x"A9" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A0" , x"CC" , x"EA" , x"F3" , x"F5" , x"F5" , x"F5" , x"EE" , x"D0" , x"D4" , x"F2" , x"F5" , x"F5" , x"DB" , x"A4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"AF" , x"EA" , x"F5" , x"F5" , x"F2" , x"B7" , x"96" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"9A" , x"CB" , x"F1" , x"F5" , x"EF" , x"BF" , x"97" , x"AE" , x"E9" , x"F5" , x"F5" , x"E3" , x"AA" , x"93" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"B0" , x"E5" , x"F5" , x"F5" , x"F0" , x"B4" , x"93" , x"92" , x"92" , x"92" , x"92" , x"92" , x"BA" , x"EC" , x"F5" , x"F5" , x"F5" , x"B4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A8" , x"E1" , x"F5" , x"F5" , x"F5" , x"D0" , x"CC" , x"EE" , x"F5" , x"F5" , x"F3" , x"D9" , x"A8" , x"93" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"AF" , x"E5" , x"F5" , x"F5" , x"EF" , x"BB" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"B4" , x"EA" , x"F5" , x"F5" , x"EC" , x"B8" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A1" , x"D3" , x"EA" , x"E6" , x"E5" , x"C9" , x"9D" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"CA" , x"F0" , x"F5" , x"F5" , x"ED" , x"B8" , x"96" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A6" , x"DB" , x"F3" , x"F5" , x"F5" , x"E3" , x"AA" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A6" , x"DC" , x"F3" , x"F5" , x"F5" , x"F0" , x"DE" , x"BA" , x"9E" , x"C1" , x"F0" , x"F5" , x"F5" , x"DB" , x"A4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"98" , x"DF" , x"F4" , x"F5" , x"F4" , x"CA" , x"9A" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A7" , x"DC" , x"F4" , x"F5" , x"E6" , x"B3" , x"94" , x"A0" , x"DC" , x"F3" , x"F5" , x"ED" , x"BE" , x"97" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"93" , x"BD" , x"ED" , x"F5" , x"F5" , x"E5" , x"AA" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"BA" , x"EC" , x"F5" , x"F5" , x"F5" , x"B4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A8" , x"E1" , x"F5" , x"F5" , x"F5" , x"CE" , x"A8" , x"D2" , x"F1" , x"F5" , x"F5" , x"F1" , x"CC" , x"9D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"AF" , x"E5" , x"F5" , x"F5" , x"EF" , x"BB" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"AF" , x"E6" , x"F5" , x"F5" , x"F2" , x"CC" , x"9C" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"95" , x"9E" , x"A2" , x"A1" , x"A1" , x"9C" , x"94" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"CA" , x"F0" , x"F5" , x"F5" , x"ED" , x"B8" , x"96" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A8" , x"DD" , x"F3" , x"F5" , x"F5" , x"DD" , x"A7" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A6" , x"DC" , x"F3" , x"F0" , x"DF" , x"C4" , x"A8" , x"97" , x"93" , x"C1" , x"F0" , x"F5" , x"F5" , x"DB" , x"A4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"94" , x"D1" , x"F1" , x"F5" , x"F4" , x"D9" , x"9D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"93" , x"B2" , x"E8" , x"F5" , x"F5" , x"D9" , x"A3" , x"93" , x"9C" , x"CF" , x"F1" , x"F5" , x"F2" , x"CA" , x"9A" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"9B" , x"CD" , x"F2" , x"F5" , x"F5" , x"D3" , x"9F" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"BA" , x"EC" , x"F5" , x"F5" , x"F5" , x"B4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A8" , x"E1" , x"F5" , x"F5" , x"F5" , x"CE" , x"9B" , x"AE" , x"E1" , x"F4" , x"F5" , x"F5" , x"EA" , x"B7" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"AF" , x"E5" , x"F5" , x"F5" , x"EF" , x"BB" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A7" , x"DD" , x"F4" , x"F5" , x"F5" , x"E8" , x"BD" , x"9A" , x"93" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"CA" , x"F0" , x"F5" , x"F5" , x"ED" , x"B8" , x"96" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"93" , x"B2" , x"E6" , x"F4" , x"F5" , x"F5" , x"D0" , x"9E" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A6" , x"D5" , x"DC" , x"C0" , x"AA" , x"99" , x"94" , x"92" , x"92" , x"C1" , x"F0" , x"F5" , x"F5" , x"DB" , x"A4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"93" , x"C2" , x"EE" , x"F5" , x"F5" , x"E4" , x"A6" , x"93" , x"92" , x"92" , x"92" , x"92" , x"92" , x"99" , x"C5" , x"EF" , x"F5" , x"F1" , x"CB" , x"9A" , x"92" , x"95" , x"BB" , x"EC" , x"F5" , x"F4" , x"D9" , x"A5" , x"93" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A5" , x"DA" , x"F3" , x"F5" , x"F1" , x"C1" , x"96" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"BA" , x"EC" , x"F5" , x"F5" , x"F5" , x"B4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A8" , x"E1" , x"F5" , x"F5" , x"F5" , x"CE" , x"9A" , x"9A" , x"C3" , x"EE" , x"F5" , x"F5" , x"F4" , x"DD" , x"A4" , x"93" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"AF" , x"E5" , x"F5" , x"F5" , x"EF" , x"BB" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"99" , x"C7" , x"F0" , x"F5" , x"F5" , x"F5" , x"E8" , x"CC" , x"B5" , x"9E" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"CA" , x"F0" , x"F5" , x"F5" , x"ED" , x"B8" , x"96" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"9D" , x"CE" , x"EF" , x"F5" , x"F5" , x"F2" , x"C1" , x"97" , x"92" , x"92" , x"92" , x"92" , x"92" , x"97" , x"A4" , x"A2" , x"96" , x"93" , x"92" , x"92" , x"92" , x"92" , x"C1" , x"F0" , x"F5" , x"F5" , x"DB" , x"A4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A8" , x"E5" , x"F5" , x"F5" , x"EC" , x"B8" , x"96" , x"92" , x"92" , x"92" , x"92" , x"92" , x"9F" , x"D7" , x"F2" , x"F5" , x"EC" , x"BA" , x"96" , x"92" , x"92" , x"AC" , x"E1" , x"F4" , x"F5" , x"E8" , x"B4" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"AD" , x"E4" , x"F4" , x"F5" , x"E8" , x"B4" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"BA" , x"EC" , x"F5" , x"F5" , x"F5" , x"B4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A8" , x"E1" , x"F5" , x"F5" , x"F5" , x"CE" , x"9A" , x"92" , x"9C" , x"D1" , x"F2" , x"F5" , x"F5" , x"F1" , x"CA" , x"9D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"AF" , x"E5" , x"F5" , x"F5" , x"EF" , x"BB" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A7" , x"DC" , x"F3" , x"F5" , x"F5" , x"F5" , x"F1" , x"EA" , x"DE" , x"CD" , x"BB" , x"A7" , x"9B" , x"98" , x"94" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"CA" , x"F0" , x"F5" , x"F5" , x"ED" , x"B8" , x"96" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"9C" , x"C7" , x"EB" , x"F5" , x"F5" , x"F5" , x"E2" , x"AF" , x"94" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"C1" , x"F0" , x"F5" , x"F5" , x"DB" , x"A4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"9F" , x"D8" , x"F2" , x"F5" , x"F0" , x"C7" , x"98" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A9" , x"E4" , x"F4" , x"F5" , x"E3" , x"A8" , x"94" , x"92" , x"92" , x"A1" , x"D5" , x"F3" , x"F5" , x"F1" , x"C3" , x"97" , x"92" , x"92" , x"92" , x"92" , x"94" , x"B8" , x"EC" , x"F5" , x"F5" , x"DD" , x"A7" , x"93" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"BA" , x"EC" , x"F5" , x"F5" , x"F5" , x"B4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A8" , x"E1" , x"F5" , x"F5" , x"F5" , x"CE" , x"9A" , x"92" , x"92" , x"AD" , x"E3" , x"F4" , x"F5" , x"F5" , x"EA" , x"BA" , x"97" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"AF" , x"E5" , x"F5" , x"F5" , x"EF" , x"BB" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"94" , x"B2" , x"DF" , x"F3" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F1" , x"EE" , x"E7" , x"DD" , x"CF" , x"BD" , x"AB" , x"A3" , x"9A" , x"93" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"CA" , x"F0" , x"F5" , x"F5" , x"ED" , x"B8" , x"96" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A1" , x"AA" , x"B3" , x"CC" , x"EC" , x"F4" , x"F5" , x"F5" , x"F1" , x"CA" , x"9B" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"C1" , x"F0" , x"F5" , x"F5" , x"DB" , x"A4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"9B" , x"CB" , x"F0" , x"F5" , x"F4" , x"D2" , x"9D" , x"92" , x"92" , x"92" , x"92" , x"93" , x"BE" , x"ED" , x"F5" , x"F4" , x"D3" , x"9C" , x"92" , x"92" , x"92" , x"97" , x"C5" , x"F0" , x"F5" , x"F5" , x"D6" , x"A1" , x"92" , x"92" , x"92" , x"92" , x"9B" , x"CC" , x"F0" , x"F5" , x"F2" , x"CC" , x"9B" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"BA" , x"EC" , x"F5" , x"F5" , x"F5" , x"B4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A8" , x"E1" , x"F5" , x"F5" , x"F5" , x"CE" , x"9A" , x"92" , x"92" , x"96" , x"BF" , x"EB" , x"F5" , x"F5" , x"F3" , x"DC" , x"AB" , x"93" , x"92" , x"92" , x"92" , x"92" , x"92" , x"AF" , x"E5" , x"F5" , x"F5" , x"EF" , x"BB" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"96" , x"B1" , x"D5" , x"EE" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F4" , x"F1" , x"ED" , x"E5" , x"DB" , x"CA" , x"B6" , x"A5" , x"97" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"CA" , x"F0" , x"F5" , x"F5" , x"F2" , x"DB" , x"CC" , x"CB" , x"CB" , x"CB" , x"CB" , x"CB" , x"CB" , x"CB" , x"CB" , x"CB" , x"D8" , x"E0" , x"E8" , x"F0" , x"F5" , x"F5" , x"F5" , x"F5" , x"DF" , x"AA" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"C1" , x"F0" , x"F5" , x"F5" , x"DB" , x"A4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"95" , x"B7" , x"EA" , x"F5" , x"F5" , x"DF" , x"AA" , x"93" , x"92" , x"92" , x"92" , x"95" , x"D0" , x"F1" , x"F5" , x"F3" , x"C3" , x"99" , x"92" , x"92" , x"92" , x"92" , x"B6" , x"EA" , x"F5" , x"F5" , x"E4" , x"AA" , x"92" , x"92" , x"92" , x"92" , x"9F" , x"D9" , x"F2" , x"F5" , x"EE" , x"C0" , x"97" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"BA" , x"EC" , x"F5" , x"F5" , x"F5" , x"B4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A8" , x"E1" , x"F5" , x"F5" , x"F5" , x"CE" , x"9A" , x"92" , x"92" , x"92" , x"A0" , x"D3" , x"F1" , x"F5" , x"F5" , x"F0" , x"CB" , x"9C" , x"92" , x"92" , x"92" , x"92" , x"92" , x"AF" , x"E5" , x"F5" , x"F5" , x"EF" , x"BB" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"96" , x"A4" , x"BE" , x"DE" , x"F1" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F3" , x"F0" , x"E9" , x"DB" , x"C3" , x"A4" , x"94" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"CA" , x"F0" , x"F5" , x"F5" , x"F5" , x"F5" , x"F4" , x"F4" , x"F4" , x"F4" , x"F4" , x"F4" , x"F4" , x"F4" , x"F4" , x"F4" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F3" , x"E0" , x"AB" , x"94" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"C1" , x"F0" , x"F5" , x"F5" , x"DB" , x"A4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A9" , x"DF" , x"F4" , x"F5" , x"EA" , x"B7" , x"94" , x"92" , x"92" , x"92" , x"A0" , x"E3" , x"F4" , x"F5" , x"EE" , x"A8" , x"93" , x"92" , x"92" , x"92" , x"92" , x"A6" , x"DF" , x"F5" , x"F5" , x"F2" , x"B5" , x"93" , x"92" , x"92" , x"92" , x"A9" , x"E6" , x"F5" , x"F5" , x"E5" , x"AB" , x"93" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"BA" , x"EC" , x"F5" , x"F5" , x"F5" , x"B4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A8" , x"E1" , x"F5" , x"F5" , x"F5" , x"CE" , x"9A" , x"92" , x"92" , x"92" , x"93" , x"AB" , x"DE" , x"F3" , x"F5" , x"F5" , x"EE" , x"BA" , x"96" , x"92" , x"92" , x"92" , x"92" , x"AF" , x"E5" , x"F5" , x"F5" , x"EF" , x"BB" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"95" , x"9F" , x"AE" , x"C9" , x"DD" , x"EA" , x"EF" , x"F2" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F4" , x"F0" , x"DF" , x"BA" , x"9B" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"CA" , x"F0" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F2" , x"E9" , x"D4" , x"AE" , x"94" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"C1" , x"F0" , x"F5" , x"F5" , x"DB" , x"A4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A0" , x"D2" , x"F2" , x"F5" , x"F0" , x"C0" , x"95" , x"92" , x"92" , x"92" , x"B5" , x"ED" , x"F5" , x"F5" , x"E0" , x"9F" , x"92" , x"92" , x"92" , x"92" , x"92" , x"95" , x"CE" , x"F3" , x"F5" , x"F5" , x"CE" , x"9B" , x"92" , x"92" , x"94" , x"BF" , x"ED" , x"F5" , x"F4" , x"D8" , x"9F" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"BA" , x"EC" , x"F5" , x"F5" , x"F5" , x"B4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A8" , x"E1" , x"F5" , x"F5" , x"F5" , x"CE" , x"9A" , x"92" , x"92" , x"92" , x"92" , x"95" , x"BB" , x"E9" , x"F5" , x"F5" , x"F5" , x"E1" , x"A8" , x"94" , x"92" , x"92" , x"92" , x"AF" , x"E5" , x"F5" , x"F5" , x"EF" , x"BB" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"94" , x"9A" , x"9F" , x"AE" , x"C1" , x"CE" , x"DB" , x"E8" , x"EF" , x"F3" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F3" , x"E7" , x"C0" , x"9D" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"CA" , x"F0" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F2" , x"ED" , x"E7" , x"DD" , x"C8" , x"B7" , x"A2" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"C1" , x"F0" , x"F5" , x"F5" , x"DB" , x"A4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"95" , x"C2" , x"EF" , x"F5" , x"F4" , x"CD" , x"9C" , x"92" , x"92" , x"92" , x"C6" , x"F1" , x"F5" , x"F5" , x"CD" , x"98" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"C0" , x"F0" , x"F5" , x"F5" , x"E1" , x"9F" , x"92" , x"92" , x"95" , x"D0" , x"F1" , x"F5" , x"F3" , x"C8" , x"9A" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"BA" , x"EC" , x"F5" , x"F5" , x"F5" , x"B4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A8" , x"E1" , x"F5" , x"F5" , x"F5" , x"CE" , x"9A" , x"92" , x"92" , x"92" , x"92" , x"92" , x"9E" , x"D2" , x"F2" , x"F5" , x"F5" , x"F2" , x"CD" , x"9E" , x"92" , x"92" , x"92" , x"AF" , x"E5" , x"F5" , x"F5" , x"EF" , x"BB" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"94" , x"97" , x"9A" , x"A3" , x"B3" , x"BE" , x"CC" , x"DF" , x"ED" , x"F4" , x"F5" , x"F5" , x"F5" , x"F4" , x"E7" , x"B8" , x"96" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"CA" , x"F0" , x"F5" , x"F5" , x"F0" , x"D0" , x"BA" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B4" , x"B2" , x"AD" , x"A5" , x"98" , x"95" , x"93" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"C1" , x"F0" , x"F5" , x"F5" , x"DB" , x"A4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"B4" , x"E8" , x"F5" , x"F5" , x"DF" , x"A7" , x"92" , x"92" , x"9B" , x"D5" , x"F4" , x"F5" , x"F1" , x"B7" , x"94" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"AD" , x"EA" , x"F5" , x"F5" , x"EE" , x"AA" , x"94" , x"92" , x"96" , x"DE" , x"F4" , x"F5" , x"EF" , x"AF" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"BA" , x"EC" , x"F5" , x"F5" , x"F5" , x"B4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A8" , x"E1" , x"F5" , x"F5" , x"F5" , x"CE" , x"9A" , x"92" , x"92" , x"92" , x"92" , x"92" , x"93" , x"A8" , x"E1" , x"F4" , x"F5" , x"F5" , x"EA" , x"BA" , x"96" , x"92" , x"92" , x"AF" , x"E5" , x"F5" , x"F5" , x"EF" , x"BB" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"93" , x"95" , x"96" , x"9A" , x"A7" , x"B4" , x"D6" , x"EE" , x"F4" , x"F5" , x"F5" , x"F4" , x"DB" , x"A2" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"CA" , x"F0" , x"F5" , x"F5" , x"ED" , x"B8" , x"96" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"C1" , x"F0" , x"F5" , x"F5" , x"DB" , x"A4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A5" , x"DD" , x"F5" , x"F5" , x"EB" , x"AF" , x"92" , x"92" , x"AD" , x"E3" , x"F5" , x"F5" , x"E5" , x"AB" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"98" , x"DC" , x"F3" , x"F5" , x"F2" , x"C0" , x"98" , x"92" , x"AC" , x"EA" , x"F5" , x"F5" , x"E4" , x"A0" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"BA" , x"EC" , x"F5" , x"F5" , x"F5" , x"B4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A8" , x"E1" , x"F5" , x"F5" , x"F5" , x"CE" , x"9A" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"94" , x"BE" , x"E9" , x"F5" , x"F5" , x"F4" , x"E0" , x"AE" , x"95" , x"92" , x"AF" , x"E5" , x"F5" , x"F5" , x"EF" , x"BB" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"93" , x"9D" , x"BB" , x"E3" , x"F4" , x"F5" , x"F5" , x"F1" , x"B9" , x"95" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"CA" , x"F0" , x"F5" , x"F5" , x"ED" , x"B8" , x"96" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"C1" , x"F0" , x"F5" , x"F5" , x"DB" , x"A4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"95" , x"CF" , x"F3" , x"F5" , x"F2" , x"BB" , x"94" , x"92" , x"BA" , x"EC" , x"F5" , x"F5" , x"D4" , x"A0" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"95" , x"CD" , x"F0" , x"F5" , x"F4" , x"CE" , x"9B" , x"92" , x"BD" , x"EF" , x"F5" , x"F5" , x"D4" , x"9B" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"BA" , x"EC" , x"F5" , x"F5" , x"F5" , x"B4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A8" , x"E1" , x"F5" , x"F5" , x"F5" , x"CE" , x"9A" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"9F" , x"CD" , x"EF" , x"F5" , x"F5" , x"F2" , x"D0" , x"9F" , x"92" , x"AF" , x"E5" , x"F5" , x"F5" , x"EF" , x"BB" , x"95" , x"92" , x"92" , x"92" , x"93" , x"A0" , x"AA" , x"AE" , x"AF" , x"AA" , x"96" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"9A" , x"C0" , x"ED" , x"F5" , x"F5" , x"F5" , x"CF" , x"9B" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"CA" , x"F0" , x"F5" , x"F5" , x"ED" , x"B8" , x"96" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"C1" , x"F0" , x"F5" , x"F5" , x"DB" , x"A4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"C0" , x"EF" , x"F5" , x"F5" , x"D0" , x"9A" , x"99" , x"CA" , x"F2" , x"F5" , x"F1" , x"C1" , x"97" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"93" , x"BA" , x"EC" , x"F5" , x"F5" , x"DC" , x"9E" , x"92" , x"CA" , x"F2" , x"F5" , x"F3" , x"BC" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"BA" , x"EC" , x"F5" , x"F5" , x"F5" , x"B4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A8" , x"E1" , x"F5" , x"F5" , x"F5" , x"CE" , x"9A" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"93" , x"AA" , x"DE" , x"F4" , x"F5" , x"F5" , x"ED" , x"BC" , x"97" , x"AF" , x"E5" , x"F5" , x"F5" , x"EF" , x"BB" , x"95" , x"92" , x"92" , x"92" , x"95" , x"C1" , x"DF" , x"E5" , x"E8" , x"D9" , x"A1" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A0" , x"DF" , x"F5" , x"F5" , x"F5" , x"D8" , x"9D" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"CA" , x"F0" , x"F5" , x"F5" , x"ED" , x"B8" , x"96" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"C1" , x"F0" , x"F5" , x"F5" , x"DB" , x"A4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"AE" , x"E9" , x"F5" , x"F5" , x"DF" , x"9F" , x"A5" , x"DA" , x"F3" , x"F5" , x"E9" , x"B6" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A6" , x"E1" , x"F4" , x"F5" , x"E8" , x"AF" , x"A1" , x"D9" , x"F5" , x"F5" , x"E9" , x"AE" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"BA" , x"EC" , x"F5" , x"F5" , x"F5" , x"B4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A8" , x"E1" , x"F5" , x"F5" , x"F5" , x"CE" , x"9A" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"97" , x"BB" , x"EA" , x"F5" , x"F5" , x"F5" , x"E4" , x"AA" , x"B1" , x"E5" , x"F5" , x"F5" , x"EF" , x"BB" , x"95" , x"92" , x"92" , x"92" , x"96" , x"C8" , x"EF" , x"F5" , x"F5" , x"E8" , x"B2" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"93" , x"D2" , x"F4" , x"F5" , x"F5" , x"DD" , x"9E" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"CA" , x"F0" , x"F5" , x"F5" , x"ED" , x"B8" , x"96" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"C1" , x"F0" , x"F5" , x"F5" , x"DB" , x"A4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"98" , x"DE" , x"F4" , x"F5" , x"EA" , x"A5" , x"AE" , x"E4" , x"F5" , x"F5" , x"DC" , x"A6" , x"93" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"9D" , x"D2" , x"F1" , x"F5" , x"ED" , x"BF" , x"B4" , x"E5" , x"F5" , x"F5" , x"DB" , x"A4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"BA" , x"EC" , x"F5" , x"F5" , x"F5" , x"B4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A8" , x"E1" , x"F5" , x"F5" , x"F5" , x"CE" , x"9A" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"97" , x"CA" , x"F1" , x"F5" , x"F5" , x"F3" , x"D1" , x"BE" , x"E6" , x"F5" , x"F5" , x"EF" , x"BB" , x"95" , x"92" , x"92" , x"92" , x"94" , x"BA" , x"EC" , x"F5" , x"F5" , x"F0" , x"C7" , x"99" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"95" , x"D3" , x"F4" , x"F5" , x"F5" , x"D9" , x"9D" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"CA" , x"F0" , x"F5" , x"F5" , x"ED" , x"B8" , x"96" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"C1" , x"F0" , x"F5" , x"F5" , x"DB" , x"A4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"94" , x"CF" , x"F0" , x"F5" , x"F2" , x"B6" , x"BE" , x"EC" , x"F5" , x"F3" , x"CE" , x"9A" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"96" , x"BF" , x"EE" , x"F5" , x"F1" , x"C7" , x"C0" , x"EC" , x"F5" , x"F4" , x"C9" , x"9A" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"BA" , x"EC" , x"F5" , x"F5" , x"F5" , x"B4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A8" , x"E1" , x"F5" , x"F5" , x"F5" , x"CE" , x"9A" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A8" , x"E0" , x"F4" , x"F5" , x"F5" , x"EB" , x"DB" , x"EB" , x"F5" , x"F5" , x"EF" , x"BB" , x"95" , x"92" , x"92" , x"92" , x"92" , x"A7" , x"E2" , x"F4" , x"F5" , x"F5" , x"DF" , x"AA" , x"93" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A5" , x"E0" , x"F5" , x"F5" , x"F5" , x"D0" , x"9B" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"CA" , x"F0" , x"F5" , x"F5" , x"ED" , x"B8" , x"96" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"C1" , x"F0" , x"F5" , x"F5" , x"DB" , x"A4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"93" , x"BD" , x"ED" , x"F5" , x"F3" , x"CF" , x"D5" , x"F0" , x"F5" , x"ED" , x"C0" , x"98" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"AE" , x"E6" , x"F5" , x"F3" , x"D4" , x"CF" , x"F0" , x"F5" , x"ED" , x"BB" , x"94" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"BA" , x"EC" , x"F5" , x"F5" , x"F5" , x"B4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A8" , x"E1" , x"F5" , x"F5" , x"F5" , x"CE" , x"9A" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"95" , x"B8" , x"E9" , x"F5" , x"F5" , x"F4" , x"F0" , x"F2" , x"F5" , x"F5" , x"EF" , x"BB" , x"95" , x"92" , x"92" , x"92" , x"92" , x"9D" , x"CF" , x"F1" , x"F5" , x"F5" , x"F0" , x"D1" , x"A0" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"99" , x"C2" , x"ED" , x"F5" , x"F5" , x"F1" , x"B9" , x"95" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"CA" , x"F0" , x"F5" , x"F5" , x"ED" , x"B8" , x"96" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"C1" , x"F0" , x"F5" , x"F5" , x"DB" , x"A4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"A7" , x"E4" , x"F5" , x"F4" , x"E0" , x"E6" , x"F3" , x"F5" , x"E6" , x"AB" , x"94" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A5" , x"DB" , x"F3" , x"F5" , x"E6" , x"E2" , x"F3" , x"F5" , x"E2" , x"AD" , x"93" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"BA" , x"EC" , x"F5" , x"F5" , x"F5" , x"B4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A8" , x"E1" , x"F5" , x"F5" , x"F5" , x"CE" , x"9A" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"9B" , x"CB" , x"F0" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"EF" , x"BB" , x"95" , x"92" , x"92" , x"92" , x"92" , x"93" , x"B1" , x"E3" , x"F5" , x"F5" , x"F5" , x"F1" , x"D5" , x"AA" , x"98" , x"93" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"94" , x"9D" , x"C1" , x"E6" , x"F5" , x"F5" , x"F4" , x"DE" , x"A5" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"CA" , x"F0" , x"F5" , x"F5" , x"ED" , x"B8" , x"96" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"C1" , x"F0" , x"F5" , x"F5" , x"DB" , x"A4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"9E" , x"D7" , x"F2" , x"F5" , x"ED" , x"F3" , x"F5" , x"F4" , x"D7" , x"9E" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"9A" , x"CB" , x"F1" , x"F5" , x"EF" , x"EE" , x"F5" , x"F3" , x"D1" , x"9D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"BA" , x"EC" , x"F5" , x"F5" , x"F5" , x"B4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A8" , x"E1" , x"F5" , x"F5" , x"F5" , x"CE" , x"9A" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"93" , x"A8" , x"D9" , x"F2" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"EF" , x"BB" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"9A" , x"C3" , x"EE" , x"F5" , x"F5" , x"F5" , x"F2" , x"E3" , x"CA" , x"AF" , x"A4" , x"9D" , x"95" , x"92" , x"92" , x"97" , x"9E" , x"A4" , x"B2" , x"D2" , x"EB" , x"F4" , x"F5" , x"F5" , x"EA" , x"BA" , x"97" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"CA" , x"F0" , x"F5" , x"F5" , x"ED" , x"B8" , x"96" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"C1" , x"F0" , x"F5" , x"F5" , x"DB" , x"A4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"99" , x"C6" , x"F0" , x"F5" , x"F4" , x"F5" , x"F5" , x"F3" , x"C4" , x"99" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"BA" , x"EC" , x"F5" , x"F4" , x"F4" , x"F5" , x"F0" , x"C5" , x"98" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"BA" , x"EC" , x"F5" , x"F5" , x"F5" , x"B4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A8" , x"E1" , x"F5" , x"F5" , x"F5" , x"CE" , x"9A" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"94" , x"B7" , x"E9" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"EF" , x"BB" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A0" , x"D1" , x"F1" , x"F5" , x"F5" , x"F5" , x"F4" , x"F0" , x"E6" , x"DA" , x"CE" , x"C2" , x"BD" , x"BD" , x"C5" , x"D1" , x"DC" , x"E9" , x"F1" , x"F5" , x"F5" , x"F5" , x"ED" , x"C9" , x"9F" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"CA" , x"F0" , x"F5" , x"F5" , x"ED" , x"B8" , x"96" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"C1" , x"F0" , x"F5" , x"F5" , x"DB" , x"A4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"94" , x"B5" , x"E9" , x"F5" , x"F5" , x"F5" , x"F5" , x"F1" , x"AE" , x"94" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"AC" , x"E3" , x"F5" , x"F5" , x"F5" , x"F5" , x"EA" , x"B5" , x"96" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"BA" , x"EC" , x"F5" , x"F5" , x"F5" , x"B4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A8" , x"E1" , x"F5" , x"F5" , x"F5" , x"CE" , x"9A" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"9B" , x"CD" , x"F1" , x"F5" , x"F5" , x"F5" , x"F5" , x"EF" , x"BB" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A5" , x"CF" , x"ED" , x"F5" , x"F5" , x"F5" , x"F5" , x"F4" , x"F3" , x"F2" , x"F0" , x"EF" , x"EF" , x"F1" , x"F3" , x"F4" , x"F5" , x"F5" , x"F5" , x"F5" , x"EF" , x"CB" , x"A2" , x"94" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"CA" , x"F0" , x"F5" , x"F5" , x"ED" , x"B8" , x"96" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"C1" , x"F0" , x"F5" , x"F5" , x"DB" , x"A4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A9" , x"DF" , x"F4" , x"F5" , x"F5" , x"F5" , x"E3" , x"A0" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"97" , x"D3" , x"F5" , x"F5" , x"F5" , x"F5" , x"DD" , x"A1" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"BA" , x"EC" , x"F5" , x"F5" , x"F5" , x"B4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A8" , x"E1" , x"F5" , x"F5" , x"F5" , x"CE" , x"9A" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"9F" , x"DB" , x"F2" , x"F5" , x"F5" , x"F5" , x"EF" , x"BB" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"9D" , x"B9" , x"DC" , x"ED" , x"F3" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F4" , x"EE" , x"DE" , x"B9" , x"9C" , x"93" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"CA" , x"F0" , x"F5" , x"F5" , x"ED" , x"B8" , x"96" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"C1" , x"F0" , x"F5" , x"F5" , x"DB" , x"A4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"9D" , x"D0" , x"F2" , x"F5" , x"F5" , x"F5" , x"D1" , x"99" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"C4" , x"F1" , x"F5" , x"F5" , x"F4" , x"CF" , x"9B" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"BA" , x"EC" , x"F5" , x"F5" , x"F5" , x"B4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A8" , x"E1" , x"F5" , x"F5" , x"F5" , x"CE" , x"9A" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"94" , x"B7" , x"E6" , x"F4" , x"F5" , x"F5" , x"EF" , x"BB" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"97" , x"A5" , x"BE" , x"D2" , x"E2" , x"E9" , x"EE" , x"F2" , x"F5" , x"F5" , x"F5" , x"F4" , x"F1" , x"ED" , x"E5" , x"D4" , x"C1" , x"A7" , x"97" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"B1" , x"C4" , x"C7" , x"C7" , x"C2" , x"A7" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"AB" , x"C4" , x"C7" , x"C7" , x"B9" , x"9D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"93" , x"AD" , x"C5" , x"C7" , x"C7" , x"C7" , x"AC" , x"94" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A8" , x"C3" , x"C7" , x"C7" , x"C6" , x"AD" , x"96" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"A8" , x"C3" , x"C7" , x"C7" , x"C7" , x"A4" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"9D" , x"BC" , x"C7" , x"C7" , x"C7" , x"B2" , x"96" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"9B" , x"B8" , x"C5" , x"C7" , x"C7" , x"C4" , x"A9" , x"94" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"93" , x"98" , x"9E" , x"AC" , x"B5" , x"BD" , x"C3" , x"C6" , x"C7" , x"C7" , x"C6" , x"C1" , x"BB" , x"B0" , x"9E" , x"97" , x"94" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"95" , x"96" , x"96" , x"96" , x"95" , x"94" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"94" , x"96" , x"96" , x"96" , x"95" , x"93" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"94" , x"96" , x"96" , x"96" , x"96" , x"94" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"94" , x"96" , x"96" , x"96" , x"96" , x"94" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"94" , x"95" , x"96" , x"96" , x"96" , x"93" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"93" , x"95" , x"96" , x"96" , x"96" , x"95" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"95" , x"96" , x"96" , x"96" , x"96" , x"94" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"94" , x"95" , x"95" , x"95" , x"96" , x"96" , x"96" , x"96" , x"96" , x"95" , x"94" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" )
);




CONSTANT P2winsR : ImageMatrix(0 TO 99, 0 TO 199) := (
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"BC" , x"C1" , x"C2" , x"C4" , x"C5" , x"C5" , x"C4" , x"C1" , x"C0" , x"BD" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"C2" , x"CB" , x"CD" , x"CD" , x"CD" , x"CD" , x"CD" , x"CD" , x"CD" , x"CD" , x"CD" , x"CD" , x"CD" , x"CD" , x"CD" , x"CD" , x"CD" , x"C9" , x"C6" , x"C3" , x"BC" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"C1" , x"CB" , x"CD" , x"CD" , x"CB" , x"C0" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BE" , x"CB" , x"CD" , x"CD" , x"CD" , x"CD" , x"C3" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BA" , x"C9" , x"CD" , x"CD" , x"CD" , x"C4" , x"B9" , x"B7" , x"B7" , x"B7" , x"BF" , x"CB" , x"CD" , x"CD" , x"CD" , x"BE" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BB" , x"C7" , x"CD" , x"CD" , x"CD" , x"CB" , x"BC" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BE" , x"C9" , x"CD" , x"CD" , x"CC" , x"C1" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BA" , x"C3" , x"CD" , x"D7" , x"DD" , x"E3" , x"E7" , x"E8" , x"E8" , x"E6" , x"E1" , x"DF" , x"D8" , x"CD" , x"C4" , x"BB" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"D1" , x"E6" , x"E9" , x"E9" , x"E9" , x"E9" , x"E9" , x"E9" , x"E9" , x"E9" , x"E9" , x"E9" , x"E9" , x"E9" , x"E9" , x"E9" , x"E9" , x"E5" , x"E4" , x"E1" , x"D8" , x"CC" , x"BE" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BA" , x"C6" , x"CD" , x"D2" , x"D6" , x"D5" , x"D5" , x"CF" , x"C9" , x"C3" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"C9" , x"E4" , x"E9" , x"E9" , x"E7" , x"CF" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"CD" , x"E6" , x"E9" , x"E9" , x"E9" , x"E9" , x"D7" , x"BD" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C4" , x"E3" , x"E9" , x"E9" , x"E8" , x"D1" , x"BA" , x"B7" , x"B7" , x"B7" , x"CA" , x"E5" , x"E9" , x"E9" , x"E9" , x"C8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C0" , x"DE" , x"E9" , x"E9" , x"E9" , x"E7" , x"D0" , x"BA" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C5" , x"E1" , x"E9" , x"E9" , x"E6" , x"CB" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"C0" , x"D1" , x"E0" , x"E9" , x"EB" , x"EC" , x"EC" , x"EE" , x"ED" , x"ED" , x"ED" , x"EC" , x"EC" , x"EB" , x"E8" , x"E2" , x"D5" , x"C4" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"D4" , x"E9" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"EE" , x"ED" , x"ED" , x"EC" , x"E8" , x"E0" , x"CC" , x"BA" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"BF" , x"D0" , x"DF" , x"E6" , x"E9" , x"EA" , x"ED" , x"ED" , x"EC" , x"EA" , x"E8" , x"E4" , x"DB" , x"C7" , x"BC" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C4" , x"E1" , x"EC" , x"ED" , x"ED" , x"D8" , x"BC" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"D8" , x"EB" , x"ED" , x"ED" , x"ED" , x"ED" , x"E3" , x"C3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"D0" , x"E9" , x"ED" , x"ED" , x"E7" , x"C9" , x"B9" , x"B7" , x"B7" , x"B7" , x"CC" , x"E8" , x"ED" , x"ED" , x"ED" , x"C9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C1" , x"E1" , x"ED" , x"ED" , x"ED" , x"ED" , x"E4" , x"C8" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C5" , x"E4" , x"EC" , x"ED" , x"E9" , x"CC" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BA" , x"C9" , x"E0" , x"EA" , x"EC" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"EB" , x"E2" , x"CC" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"D4" , x"E9" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"EC" , x"E8" , x"CE" , x"BC" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B9" , x"C6" , x"DA" , x"E8" , x"EC" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"EC" , x"E6" , x"D3" , x"BE" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BE" , x"DA" , x"EB" , x"ED" , x"ED" , x"E0" , x"C0" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BC" , x"E2" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"E9" , x"C9" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"D9" , x"EB" , x"ED" , x"ED" , x"E0" , x"BF" , x"B7" , x"B7" , x"B7" , x"B7" , x"CC" , x"E8" , x"ED" , x"ED" , x"ED" , x"C9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C1" , x"E1" , x"ED" , x"ED" , x"ED" , x"ED" , x"EB" , x"DC" , x"C1" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C5" , x"E4" , x"EC" , x"ED" , x"E9" , x"CC" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C8" , x"E3" , x"EC" , x"ED" , x"ED" , x"ED" , x"EA" , x"E8" , x"E3" , x"DE" , x"DD" , x"DD" , x"DF" , x"E3" , x"E6" , x"EB" , x"ED" , x"ED" , x"ED" , x"ED" , x"E5" , x"CD" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"D4" , x"E9" , x"ED" , x"ED" , x"EA" , x"DE" , x"D5" , x"D5" , x"D5" , x"D5" , x"D5" , x"D5" , x"D5" , x"D5" , x"D5" , x"D5" , x"D6" , x"DD" , x"E3" , x"EA" , x"ED" , x"ED" , x"ED" , x"ED" , x"E3" , x"C7" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"C7" , x"DF" , x"EB" , x"ED" , x"ED" , x"ED" , x"EC" , x"E8" , x"E3" , x"E3" , x"E6" , x"EB" , x"EC" , x"ED" , x"ED" , x"EC" , x"E8" , x"D5" , x"BE" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"D1" , x"EA" , x"ED" , x"ED" , x"E6" , x"C6" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C7" , x"E7" , x"ED" , x"ED" , x"EB" , x"EC" , x"ED" , x"ED" , x"D5" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BB" , x"E1" , x"EC" , x"ED" , x"ED" , x"D6" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"CC" , x"E8" , x"ED" , x"ED" , x"ED" , x"C9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C1" , x"E1" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"E9" , x"D2" , x"BC" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C5" , x"E4" , x"EC" , x"ED" , x"E9" , x"CC" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C0" , x"DD" , x"EB" , x"ED" , x"ED" , x"EC" , x"E1" , x"D3" , x"CC" , x"C5" , x"BE" , x"BC" , x"BC" , x"BF" , x"C5" , x"CA" , x"D5" , x"E4" , x"EC" , x"ED" , x"ED" , x"EC" , x"E1" , x"C6" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"D4" , x"E9" , x"ED" , x"ED" , x"E8" , x"CC" , x"BB" , x"BA" , x"BA" , x"BA" , x"BA" , x"BA" , x"BA" , x"BA" , x"BA" , x"BA" , x"BA" , x"BF" , x"C4" , x"D2" , x"E7" , x"ED" , x"ED" , x"ED" , x"EB" , x"D9" , x"BF" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"C0" , x"DC" , x"EA" , x"ED" , x"ED" , x"EB" , x"E4" , x"D2" , x"C8" , x"C5" , x"C5" , x"C6" , x"CC" , x"DB" , x"E9" , x"ED" , x"ED" , x"ED" , x"E8" , x"D0" , x"BA" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B6" , x"CA" , x"E6" , x"ED" , x"ED" , x"EC" , x"CD" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"D1" , x"EA" , x"ED" , x"ED" , x"E1" , x"E9" , x"ED" , x"ED" , x"DF" , x"BD" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C2" , x"E5" , x"ED" , x"ED" , x"EB" , x"CE" , x"BA" , x"B7" , x"B7" , x"B7" , x"B7" , x"CC" , x"E8" , x"ED" , x"ED" , x"ED" , x"C9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C1" , x"E1" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"E5" , x"C7" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C5" , x"E4" , x"EC" , x"ED" , x"E9" , x"CC" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B9" , x"CE" , x"E7" , x"ED" , x"ED" , x"EC" , x"DB" , x"C6" , x"BA" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"B9" , x"BC" , x"C7" , x"DF" , x"EC" , x"ED" , x"ED" , x"EA" , x"D7" , x"BD" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"D4" , x"E9" , x"ED" , x"ED" , x"E8" , x"CA" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B9" , x"CC" , x"E4" , x"EC" , x"ED" , x"ED" , x"E7" , x"CB" , x"B9" , x"B7" , x"B7" , x"B7" , x"B8" , x"D4" , x"E9" , x"ED" , x"ED" , x"E9" , x"DA" , x"C3" , x"BA" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"BC" , x"CB" , x"E2" , x"EC" , x"ED" , x"ED" , x"E7" , x"C6" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C1" , x"E0" , x"ED" , x"ED" , x"ED" , x"D7" , x"BA" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BD" , x"DC" , x"EC" , x"ED" , x"E8" , x"CF" , x"E5" , x"ED" , x"ED" , x"EA" , x"C3" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"CC" , x"E9" , x"ED" , x"ED" , x"E7" , x"C2" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"CC" , x"E8" , x"ED" , x"ED" , x"ED" , x"C9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C1" , x"E1" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"DE" , x"C0" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C5" , x"E4" , x"EC" , x"ED" , x"E9" , x"CC" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C0" , x"DD" , x"ED" , x"ED" , x"EC" , x"E0" , x"C2" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"C4" , x"DE" , x"EB" , x"ED" , x"ED" , x"E4" , x"C9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"D4" , x"E9" , x"ED" , x"ED" , x"E8" , x"CA" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BB" , x"D3" , x"E9" , x"ED" , x"ED" , x"EB" , x"D3" , x"BB" , x"B7" , x"B7" , x"B7" , x"BE" , x"E2" , x"EC" , x"ED" , x"ED" , x"DC" , x"C2" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BA" , x"CD" , x"E8" , x"ED" , x"ED" , x"EC" , x"D3" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"D8" , x"EC" , x"ED" , x"ED" , x"DE" , x"BD" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C4" , x"E2" , x"ED" , x"ED" , x"E1" , x"C5" , x"DC" , x"EB" , x"ED" , x"EC" , x"CF" , x"BA" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"D6" , x"EC" , x"ED" , x"ED" , x"DE" , x"BD" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"CC" , x"E8" , x"ED" , x"ED" , x"ED" , x"C9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C1" , x"E1" , x"ED" , x"ED" , x"ED" , x"EB" , x"EC" , x"ED" , x"ED" , x"EA" , x"D2" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C5" , x"E4" , x"EC" , x"ED" , x"E9" , x"CC" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C5" , x"E2" , x"EC" , x"ED" , x"EA" , x"D0" , x"BA" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B9" , x"CF" , x"E8" , x"EE" , x"ED" , x"EB" , x"D0" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"D4" , x"E9" , x"ED" , x"ED" , x"E8" , x"CA" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C6" , x"E4" , x"EC" , x"ED" , x"ED" , x"DB" , x"BF" , x"B7" , x"B7" , x"B7" , x"CA" , x"E8" , x"ED" , x"ED" , x"EA" , x"C9" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BB" , x"DD" , x"EB" , x"ED" , x"ED" , x"DE" , x"BD" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"D0" , x"E9" , x"ED" , x"ED" , x"E7" , x"C0" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"CB" , x"E7" , x"ED" , x"EC" , x"D8" , x"BD" , x"D2" , x"E9" , x"ED" , x"EC" , x"DA" , x"BC" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BD" , x"DE" , x"EE" , x"ED" , x"ED" , x"D5" , x"BA" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"CC" , x"E8" , x"ED" , x"ED" , x"ED" , x"C9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C1" , x"E1" , x"ED" , x"ED" , x"ED" , x"E0" , x"E6" , x"EC" , x"ED" , x"ED" , x"E4" , x"CA" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C5" , x"E4" , x"EC" , x"ED" , x"E9" , x"CC" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C9" , x"E6" , x"ED" , x"ED" , x"E7" , x"CA" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C4" , x"E0" , x"ED" , x"ED" , x"ED" , x"D7" , x"BC" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"D4" , x"E9" , x"ED" , x"ED" , x"E8" , x"CA" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C1" , x"DF" , x"ED" , x"ED" , x"ED" , x"DF" , x"C2" , x"B7" , x"B7" , x"B7" , x"D4" , x"EB" , x"ED" , x"ED" , x"E1" , x"BF" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"D3" , x"E9" , x"ED" , x"ED" , x"E3" , x"BF" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C5" , x"E6" , x"ED" , x"ED" , x"EC" , x"C9" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BB" , x"D5" , x"EB" , x"ED" , x"E9" , x"CE" , x"B9" , x"C4" , x"E6" , x"ED" , x"ED" , x"E3" , x"C3" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C5" , x"E4" , x"ED" , x"ED" , x"EA" , x"CA" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"CC" , x"E8" , x"ED" , x"ED" , x"ED" , x"C9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C1" , x"E1" , x"ED" , x"ED" , x"ED" , x"D6" , x"D4" , x"E9" , x"ED" , x"ED" , x"EC" , x"DD" , x"C1" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C5" , x"E4" , x"EC" , x"ED" , x"E9" , x"CC" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C9" , x"E7" , x"ED" , x"ED" , x"E7" , x"CA" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BE" , x"D9" , x"E7" , x"E5" , x"E4" , x"D3" , x"BC" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"D4" , x"E9" , x"ED" , x"ED" , x"E8" , x"CA" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C1" , x"DD" , x"EC" , x"ED" , x"ED" , x"E2" , x"C3" , x"B7" , x"B7" , x"BA" , x"D8" , x"E9" , x"EA" , x"EB" , x"D9" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"CD" , x"E9" , x"ED" , x"ED" , x"E6" , x"C5" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BA" , x"E1" , x"EC" , x"ED" , x"EC" , x"D3" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C1" , x"DF" , x"EC" , x"ED" , x"E4" , x"C7" , x"B7" , x"BE" , x"DD" , x"EC" , x"ED" , x"E8" , x"CC" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"CD" , x"E8" , x"ED" , x"ED" , x"E3" , x"C4" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"CC" , x"E8" , x"ED" , x"ED" , x"ED" , x"C9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C1" , x"E1" , x"ED" , x"ED" , x"ED" , x"D5" , x"C2" , x"D9" , x"EB" , x"ED" , x"ED" , x"EA" , x"D4" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C5" , x"E4" , x"EC" , x"ED" , x"E9" , x"CC" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C6" , x"E4" , x"ED" , x"ED" , x"EB" , x"D6" , x"BC" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BD" , x"C0" , x"BE" , x"BE" , x"BC" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"D4" , x"E9" , x"ED" , x"ED" , x"E8" , x"CA" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C1" , x"DE" , x"ED" , x"ED" , x"ED" , x"DF" , x"C1" , x"B7" , x"B7" , x"BA" , x"C7" , x"D0" , x"D3" , x"D5" , x"CB" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"D0" , x"E8" , x"ED" , x"ED" , x"E5" , x"C2" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"D8" , x"EB" , x"ED" , x"EC" , x"DB" , x"BD" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"C8" , x"E5" , x"ED" , x"ED" , x"DD" , x"C0" , x"B8" , x"BB" , x"D6" , x"EB" , x"ED" , x"EA" , x"D5" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BB" , x"D5" , x"EB" , x"ED" , x"ED" , x"D9" , x"BD" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"CC" , x"E8" , x"ED" , x"ED" , x"ED" , x"C9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C1" , x"E1" , x"ED" , x"ED" , x"ED" , x"D5" , x"BC" , x"C6" , x"E1" , x"ED" , x"ED" , x"ED" , x"E6" , x"CA" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C5" , x"E4" , x"EC" , x"ED" , x"E9" , x"CC" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C2" , x"DE" , x"EC" , x"ED" , x"ED" , x"E5" , x"CC" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"D4" , x"E9" , x"ED" , x"ED" , x"E8" , x"CA" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C6" , x"E3" , x"EC" , x"ED" , x"ED" , x"D8" , x"BD" , x"B7" , x"B7" , x"B8" , x"B9" , x"BA" , x"BA" , x"BA" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"D7" , x"EB" , x"ED" , x"ED" , x"E2" , x"BE" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"CF" , x"E8" , x"ED" , x"ED" , x"E3" , x"C1" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BA" , x"D1" , x"E9" , x"ED" , x"EB" , x"D4" , x"BB" , x"B7" , x"B9" , x"CC" , x"E7" , x"ED" , x"EC" , x"DD" , x"C0" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C0" , x"DD" , x"EC" , x"ED" , x"EB" , x"CF" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"CC" , x"E8" , x"ED" , x"ED" , x"ED" , x"C9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C1" , x"E1" , x"ED" , x"ED" , x"ED" , x"D5" , x"BB" , x"BB" , x"D1" , x"E8" , x"ED" , x"ED" , x"ED" , x"DD" , x"C0" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C5" , x"E4" , x"EC" , x"ED" , x"E9" , x"CC" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BA" , x"D3" , x"E9" , x"ED" , x"ED" , x"EC" , x"E5" , x"D5" , x"C8" , x"BD" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"D4" , x"E9" , x"ED" , x"ED" , x"E8" , x"CA" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BC" , x"D6" , x"EA" , x"ED" , x"ED" , x"EB" , x"D1" , x"BA" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C1" , x"E3" , x"ED" , x"ED" , x"EC" , x"D8" , x"BC" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B6" , x"C3" , x"E3" , x"EC" , x"ED" , x"E7" , x"CB" , x"BA" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BD" , x"DB" , x"EB" , x"ED" , x"E8" , x"CB" , x"B9" , x"B7" , x"B7" , x"C4" , x"E1" , x"ED" , x"ED" , x"E4" , x"C8" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C5" , x"E3" , x"EC" , x"ED" , x"E4" , x"C8" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"CC" , x"E8" , x"ED" , x"ED" , x"ED" , x"C9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C1" , x"E1" , x"ED" , x"ED" , x"ED" , x"D5" , x"BB" , x"B7" , x"BC" , x"D8" , x"EC" , x"ED" , x"ED" , x"EA" , x"D4" , x"BD" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C5" , x"E4" , x"EC" , x"ED" , x"E9" , x"CC" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C2" , x"DF" , x"EC" , x"ED" , x"ED" , x"ED" , x"EB" , x"E6" , x"DF" , x"D6" , x"CB" , x"C2" , x"BC" , x"BA" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"D4" , x"E9" , x"ED" , x"ED" , x"E8" , x"CA" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BC" , x"D2" , x"E7" , x"ED" , x"ED" , x"ED" , x"E3" , x"C6" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BB" , x"D5" , x"EB" , x"ED" , x"ED" , x"EA" , x"C9" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BD" , x"DC" , x"EC" , x"ED" , x"EA" , x"D3" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C2" , x"E2" , x"EC" , x"ED" , x"E2" , x"C2" , x"B8" , x"B7" , x"B7" , x"BD" , x"D9" , x"EB" , x"ED" , x"EA" , x"D1" , x"BA" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"CB" , x"E8" , x"ED" , x"ED" , x"DF" , x"C1" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"CC" , x"E8" , x"ED" , x"ED" , x"ED" , x"C9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C1" , x"E1" , x"ED" , x"ED" , x"ED" , x"D5" , x"BB" , x"B7" , x"B7" , x"C4" , x"E3" , x"ED" , x"ED" , x"ED" , x"E5" , x"CB" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C5" , x"E4" , x"EC" , x"ED" , x"E9" , x"CC" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"C7" , x"E0" , x"EB" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"EB" , x"E8" , x"E4" , x"DE" , x"D6" , x"CD" , x"C5" , x"BF" , x"BB" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"D4" , x"E9" , x"ED" , x"ED" , x"E8" , x"CA" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BE" , x"C3" , x"C8" , x"D5" , x"E7" , x"EC" , x"ED" , x"ED" , x"EB" , x"D5" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BA" , x"CC" , x"E5" , x"ED" , x"ED" , x"EC" , x"DB" , x"BD" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BB" , x"D3" , x"EA" , x"ED" , x"EC" , x"DA" , x"BD" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"CD" , x"E7" , x"ED" , x"ED" , x"D8" , x"BC" , x"B7" , x"B7" , x"B7" , x"B9" , x"D2" , x"EB" , x"ED" , x"ED" , x"DB" , x"BE" , x"B7" , x"B7" , x"B7" , x"B7" , x"BB" , x"D5" , x"EA" , x"ED" , x"EB" , x"D6" , x"BC" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"CC" , x"E8" , x"ED" , x"ED" , x"ED" , x"C9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C1" , x"E1" , x"ED" , x"ED" , x"ED" , x"D5" , x"BB" , x"B7" , x"B7" , x"B9" , x"CE" , x"E8" , x"ED" , x"ED" , x"EC" , x"DE" , x"C3" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C5" , x"E4" , x"EC" , x"ED" , x"E9" , x"CC" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BA" , x"C7" , x"DA" , x"E8" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"EC" , x"EB" , x"E9" , x"E5" , x"DE" , x"D5" , x"CB" , x"C1" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"D4" , x"E9" , x"ED" , x"ED" , x"EB" , x"DE" , x"D7" , x"D6" , x"D6" , x"D6" , x"D6" , x"D6" , x"D6" , x"D6" , x"D6" , x"D6" , x"DB" , x"E1" , x"E6" , x"EA" , x"ED" , x"ED" , x"ED" , x"ED" , x"DF" , x"C3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B9" , x"C8" , x"E1" , x"EC" , x"ED" , x"ED" , x"E5" , x"CA" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"CB" , x"E7" , x"ED" , x"ED" , x"E0" , x"C2" , x"B8" , x"B7" , x"B7" , x"B7" , x"B8" , x"D8" , x"EB" , x"ED" , x"EC" , x"CF" , x"BA" , x"B7" , x"B7" , x"B7" , x"B6" , x"CA" , x"E6" , x"ED" , x"ED" , x"E4" , x"C3" , x"B7" , x"B7" , x"B7" , x"B7" , x"BE" , x"DD" , x"EB" , x"ED" , x"E8" , x"CE" , x"BA" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"CC" , x"E8" , x"ED" , x"ED" , x"ED" , x"C9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C1" , x"E1" , x"ED" , x"ED" , x"ED" , x"D5" , x"BB" , x"B7" , x"B7" , x"B7" , x"BE" , x"D9" , x"EB" , x"ED" , x"ED" , x"EA" , x"D5" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C5" , x"E4" , x"EC" , x"ED" , x"E9" , x"CC" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"BF" , x"CD" , x"DE" , x"EA" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"EC" , x"EB" , x"EB" , x"E6" , x"DD" , x"D0" , x"C0" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"D4" , x"E9" , x"ED" , x"ED" , x"ED" , x"ED" , x"EC" , x"EC" , x"EC" , x"EC" , x"EC" , x"EC" , x"EC" , x"EC" , x"EC" , x"EC" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"EC" , x"E0" , x"C3" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"CA" , x"E3" , x"EC" , x"ED" , x"ED" , x"E8" , x"CF" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C3" , x"E1" , x"EC" , x"ED" , x"E6" , x"CA" , x"B8" , x"B7" , x"B7" , x"B7" , x"BC" , x"E3" , x"EC" , x"ED" , x"E8" , x"C3" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C0" , x"DF" , x"ED" , x"ED" , x"EB" , x"CA" , x"B8" , x"B7" , x"B7" , x"B6" , x"C2" , x"E5" , x"ED" , x"ED" , x"E4" , x"C3" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"CC" , x"E8" , x"ED" , x"ED" , x"ED" , x"C9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C1" , x"E1" , x"ED" , x"ED" , x"ED" , x"D5" , x"BB" , x"B7" , x"B7" , x"B7" , x"B8" , x"C4" , x"DF" , x"ED" , x"ED" , x"ED" , x"E9" , x"CC" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"C5" , x"E4" , x"EC" , x"ED" , x"E9" , x"CC" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"BE" , x"C5" , x"D2" , x"DF" , x"E6" , x"E9" , x"EC" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"EC" , x"EA" , x"E0" , x"CC" , x"BC" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"D4" , x"E9" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"EB" , x"E5" , x"D9" , x"C5" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BA" , x"C9" , x"E3" , x"EB" , x"ED" , x"ED" , x"E9" , x"D5" , x"BE" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BD" , x"D9" , x"EB" , x"ED" , x"EA" , x"CF" , x"B9" , x"B7" , x"B7" , x"B7" , x"C7" , x"E7" , x"ED" , x"ED" , x"DF" , x"BD" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"D7" , x"EC" , x"ED" , x"ED" , x"D6" , x"BA" , x"B7" , x"B7" , x"B7" , x"CD" , x"E8" , x"ED" , x"EC" , x"DC" , x"BD" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"CC" , x"E8" , x"ED" , x"ED" , x"ED" , x"C9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C1" , x"E1" , x"ED" , x"ED" , x"ED" , x"D5" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"CC" , x"E7" , x"ED" , x"ED" , x"ED" , x"E1" , x"C2" , x"B8" , x"B7" , x"B7" , x"B7" , x"C5" , x"E4" , x"EC" , x"ED" , x"E9" , x"CC" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BA" , x"BD" , x"C5" , x"CF" , x"D7" , x"DE" , x"E4" , x"E9" , x"EC" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"EC" , x"E4" , x"CF" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"D4" , x"E9" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"EB" , x"E7" , x"E4" , x"DE" , x"D3" , x"CB" , x"BF" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BB" , x"CD" , x"E3" , x"EC" , x"ED" , x"ED" , x"EA" , x"D4" , x"BF" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"D0" , x"E9" , x"ED" , x"EC" , x"D6" , x"BC" , x"B7" , x"B7" , x"B7" , x"D1" , x"EA" , x"ED" , x"ED" , x"D5" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"CE" , x"E9" , x"ED" , x"ED" , x"E0" , x"BE" , x"B7" , x"B7" , x"B9" , x"D6" , x"EA" , x"ED" , x"EC" , x"D3" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"CC" , x"E8" , x"ED" , x"ED" , x"ED" , x"C9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C1" , x"E1" , x"ED" , x"ED" , x"ED" , x"D5" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BE" , x"D8" , x"EB" , x"ED" , x"ED" , x"EB" , x"D5" , x"BC" , x"B7" , x"B7" , x"B7" , x"C5" , x"E4" , x"EC" , x"ED" , x"E9" , x"CC" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"BA" , x"BB" , x"C0" , x"C8" , x"CE" , x"D6" , x"DF" , x"E8" , x"EC" , x"ED" , x"ED" , x"ED" , x"EC" , x"E4" , x"CA" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"D4" , x"E9" , x"ED" , x"ED" , x"E9" , x"D7" , x"CC" , x"CB" , x"CB" , x"CB" , x"CB" , x"CB" , x"CB" , x"CB" , x"CB" , x"CB" , x"CA" , x"C8" , x"C4" , x"C0" , x"BA" , x"B9" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BC" , x"D1" , x"E5" , x"EC" , x"ED" , x"ED" , x"EA" , x"D7" , x"BD" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B6" , x"C7" , x"E4" , x"ED" , x"ED" , x"DF" , x"C2" , x"B7" , x"B7" , x"BB" , x"DB" , x"EC" , x"ED" , x"EA" , x"CB" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C4" , x"E6" , x"ED" , x"ED" , x"E8" , x"C2" , x"B8" , x"B7" , x"B9" , x"E0" , x"EC" , x"ED" , x"E9" , x"C6" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"CC" , x"E8" , x"ED" , x"ED" , x"ED" , x"C9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C1" , x"E1" , x"ED" , x"ED" , x"ED" , x"D5" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"C2" , x"E1" , x"EC" , x"ED" , x"EE" , x"E7" , x"CC" , x"B9" , x"B7" , x"B7" , x"C5" , x"E4" , x"EC" , x"ED" , x"E9" , x"CC" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"B8" , x"B9" , x"BB" , x"C2" , x"C9" , x"DA" , x"E8" , x"ED" , x"ED" , x"ED" , x"EC" , x"DD" , x"BF" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"D4" , x"E9" , x"ED" , x"ED" , x"E8" , x"CA" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B9" , x"C1" , x"DA" , x"E9" , x"EC" , x"ED" , x"EC" , x"E5" , x"CD" , x"BD" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BF" , x"DF" , x"ED" , x"ED" , x"E7" , x"C7" , x"B7" , x"B7" , x"C4" , x"E2" , x"ED" , x"ED" , x"E3" , x"C4" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BB" , x"DE" , x"EC" , x"ED" , x"EB" , x"CF" , x"BA" , x"B7" , x"C3" , x"E6" , x"ED" , x"ED" , x"E2" , x"BF" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"CC" , x"E8" , x"ED" , x"ED" , x"ED" , x"C9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C1" , x"E1" , x"ED" , x"ED" , x"ED" , x"D5" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"CE" , x"E7" , x"ED" , x"ED" , x"ED" , x"E0" , x"C5" , x"B7" , x"B7" , x"C5" , x"E4" , x"EC" , x"ED" , x"E9" , x"CC" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"BD" , x"CC" , x"E1" , x"EC" , x"ED" , x"ED" , x"EA" , x"CB" , x"B8" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"D4" , x"E9" , x"ED" , x"ED" , x"E8" , x"CA" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BA" , x"C7" , x"DD" , x"EB" , x"ED" , x"ED" , x"ED" , x"E3" , x"CD" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"D7" , x"ED" , x"ED" , x"EC" , x"CE" , x"B8" , x"B7" , x"CC" , x"E8" , x"ED" , x"ED" , x"DA" , x"BD" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"D5" , x"EA" , x"ED" , x"ED" , x"D6" , x"BC" , x"B7" , x"CC" , x"E8" , x"ED" , x"ED" , x"D9" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"CC" , x"E8" , x"ED" , x"ED" , x"ED" , x"C9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C1" , x"E1" , x"ED" , x"ED" , x"ED" , x"D5" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BD" , x"D6" , x"EA" , x"ED" , x"ED" , x"EB" , x"D8" , x"BD" , x"B7" , x"C5" , x"E4" , x"EC" , x"ED" , x"E9" , x"CC" , x"B9" , x"B7" , x"B7" , x"B7" , x"B8" , x"BE" , x"C3" , x"C5" , x"C7" , x"C3" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BA" , x"D0" , x"E8" , x"ED" , x"ED" , x"ED" , x"D6" , x"BB" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"D4" , x"E9" , x"ED" , x"ED" , x"E8" , x"CA" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BA" , x"CD" , x"E1" , x"EC" , x"ED" , x"ED" , x"EC" , x"E0" , x"C9" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"CE" , x"E9" , x"ED" , x"ED" , x"D6" , x"BB" , x"BA" , x"D5" , x"EB" , x"ED" , x"EA" , x"D0" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"CB" , x"E8" , x"ED" , x"ED" , x"DD" , x"BE" , x"B7" , x"D4" , x"EC" , x"ED" , x"EC" , x"CE" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"CC" , x"E8" , x"ED" , x"ED" , x"ED" , x"C9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C1" , x"E1" , x"ED" , x"ED" , x"ED" , x"D5" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"C4" , x"E1" , x"ED" , x"ED" , x"ED" , x"E8" , x"CC" , x"BA" , x"C5" , x"E4" , x"EC" , x"ED" , x"E9" , x"CC" , x"B9" , x"B7" , x"B7" , x"B7" , x"B9" , x"CF" , x"DF" , x"E3" , x"E5" , x"DC" , x"BE" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BE" , x"E0" , x"ED" , x"ED" , x"ED" , x"DB" , x"BC" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"D4" , x"E9" , x"ED" , x"ED" , x"E8" , x"CA" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BA" , x"CF" , x"E5" , x"EC" , x"ED" , x"ED" , x"EA" , x"DC" , x"C5" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C5" , x"E6" , x"ED" , x"ED" , x"DF" , x"BE" , x"C0" , x"DC" , x"EC" , x"ED" , x"E5" , x"C8" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C1" , x"E1" , x"EC" , x"ED" , x"E5" , x"C5" , x"BD" , x"DD" , x"ED" , x"ED" , x"E6" , x"C5" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"CC" , x"E8" , x"ED" , x"ED" , x"ED" , x"C9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C1" , x"E1" , x"ED" , x"ED" , x"ED" , x"D5" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B9" , x"CC" , x"E6" , x"EE" , x"ED" , x"ED" , x"E2" , x"C2" , x"C6" , x"E4" , x"EC" , x"ED" , x"E9" , x"CC" , x"B9" , x"B7" , x"B7" , x"B7" , x"B8" , x"D3" , x"E9" , x"EC" , x"ED" , x"E6" , x"C7" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"D9" , x"ED" , x"ED" , x"ED" , x"DF" , x"BE" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"D4" , x"E9" , x"ED" , x"ED" , x"E8" , x"CA" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"BE" , x"D4" , x"E8" , x"EC" , x"ED" , x"ED" , x"E7" , x"D4" , x"C0" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B9" , x"DF" , x"EC" , x"ED" , x"E7" , x"C0" , x"C5" , x"E3" , x"EC" , x"ED" , x"DE" , x"C1" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BD" , x"D8" , x"EB" , x"ED" , x"E9" , x"CD" , x"C8" , x"E4" , x"ED" , x"ED" , x"DD" , x"BF" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"CC" , x"E8" , x"ED" , x"ED" , x"ED" , x"C9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C1" , x"E1" , x"ED" , x"ED" , x"ED" , x"D5" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BA" , x"D5" , x"EB" , x"ED" , x"ED" , x"EC" , x"D9" , x"CD" , x"E4" , x"EC" , x"ED" , x"E9" , x"CC" , x"B9" , x"B7" , x"B7" , x"B7" , x"B8" , x"CA" , x"E7" , x"ED" , x"ED" , x"E9" , x"D2" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B9" , x"DA" , x"ED" , x"ED" , x"ED" , x"DB" , x"BC" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"D4" , x"E9" , x"ED" , x"ED" , x"E8" , x"CA" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BE" , x"D4" , x"E7" , x"ED" , x"ED" , x"ED" , x"E6" , x"CF" , x"BC" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"D7" , x"EA" , x"ED" , x"EC" , x"C9" , x"CD" , x"E8" , x"ED" , x"EB" , x"D5" , x"BC" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BA" , x"CF" , x"E8" , x"ED" , x"EA" , x"D2" , x"CF" , x"E6" , x"ED" , x"EC" , x"D5" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"CC" , x"E8" , x"ED" , x"ED" , x"ED" , x"C9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C1" , x"E1" , x"ED" , x"ED" , x"ED" , x"D5" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C2" , x"E0" , x"EC" , x"ED" , x"ED" , x"E7" , x"DE" , x"E7" , x"ED" , x"ED" , x"E9" , x"CC" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"C2" , x"E3" , x"EC" , x"ED" , x"EC" , x"DF" , x"C4" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C0" , x"E1" , x"ED" , x"ED" , x"ED" , x"D6" , x"BB" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"D4" , x"E9" , x"ED" , x"ED" , x"E8" , x"CA" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BA" , x"D0" , x"E6" , x"EC" , x"ED" , x"EC" , x"E3" , x"CD" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"CD" , x"E8" , x"ED" , x"ED" , x"D5" , x"D9" , x"EA" , x"ED" , x"E9" , x"CD" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C6" , x"E4" , x"ED" , x"EC" , x"DA" , x"D7" , x"E9" , x"ED" , x"E7" , x"CD" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"CC" , x"E8" , x"ED" , x"ED" , x"ED" , x"C9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C1" , x"E1" , x"ED" , x"ED" , x"ED" , x"D5" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B9" , x"CC" , x"E6" , x"ED" , x"ED" , x"ED" , x"EA" , x"EB" , x"ED" , x"ED" , x"E9" , x"CC" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"BD" , x"D7" , x"EA" , x"ED" , x"ED" , x"EA" , x"D9" , x"BE" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BB" , x"CF" , x"E8" , x"ED" , x"ED" , x"EA" , x"CB" , x"B8" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"D4" , x"E9" , x"ED" , x"ED" , x"E8" , x"CA" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"CD" , x"E5" , x"EC" , x"ED" , x"ED" , x"E0" , x"C8" , x"BA" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C2" , x"E4" , x"EC" , x"EC" , x"DF" , x"E3" , x"EB" , x"ED" , x"E3" , x"C3" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C0" , x"DC" , x"ED" , x"ED" , x"E4" , x"E1" , x"EC" , x"ED" , x"E1" , x"C4" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"CC" , x"E8" , x"ED" , x"ED" , x"ED" , x"C9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C1" , x"E1" , x"ED" , x"ED" , x"ED" , x"D5" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BC" , x"D5" , x"E9" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"E9" , x"CC" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"C7" , x"E2" , x"EC" , x"ED" , x"ED" , x"E9" , x"DA" , x"C3" , x"BA" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"BC" , x"CE" , x"E4" , x"EC" , x"ED" , x"EC" , x"DF" , x"C0" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"D4" , x"E9" , x"ED" , x"ED" , x"E8" , x"CA" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C1" , x"E2" , x"EC" , x"ED" , x"ED" , x"E2" , x"C8" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BC" , x"DB" , x"EB" , x"ED" , x"E7" , x"EB" , x"ED" , x"EC" , x"DC" , x"BD" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BB" , x"D5" , x"EB" , x"ED" , x"E9" , x"E9" , x"ED" , x"EC" , x"D9" , x"BC" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"CC" , x"E8" , x"ED" , x"ED" , x"ED" , x"C9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C1" , x"E1" , x"ED" , x"ED" , x"ED" , x"D5" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"C1" , x"DD" , x"EB" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"E9" , x"CC" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BA" , x"D0" , x"E8" , x"ED" , x"ED" , x"ED" , x"EB" , x"E3" , x"D4" , x"C6" , x"BF" , x"BB" , x"B9" , x"B7" , x"B6" , x"B9" , x"BC" , x"C0" , x"C7" , x"D8" , x"E7" , x"EC" , x"ED" , x"ED" , x"E6" , x"CC" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"D4" , x"E9" , x"ED" , x"ED" , x"E8" , x"CA" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B9" , x"D2" , x"EA" , x"ED" , x"ED" , x"ED" , x"E1" , x"D2" , x"CE" , x"CD" , x"CD" , x"CD" , x"CD" , x"CD" , x"CD" , x"CD" , x"CD" , x"CD" , x"CD" , x"CD" , x"CD" , x"CD" , x"CB" , x"BF" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B9" , x"D2" , x"EA" , x"ED" , x"EC" , x"EE" , x"ED" , x"EC" , x"D0" , x"BA" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"CC" , x"E8" , x"ED" , x"EC" , x"EC" , x"ED" , x"E9" , x"D1" , x"BA" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"CC" , x"E8" , x"ED" , x"ED" , x"ED" , x"C9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C1" , x"E1" , x"ED" , x"ED" , x"ED" , x"D5" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"CA" , x"E6" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"E9" , x"CC" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BD" , x"D8" , x"EB" , x"ED" , x"ED" , x"ED" , x"EC" , x"EA" , x"E4" , x"DC" , x"D7" , x"D1" , x"CF" , x"CE" , x"D1" , x"D6" , x"DD" , x"E5" , x"EB" , x"ED" , x"ED" , x"ED" , x"E8" , x"D3" , x"BE" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"D4" , x"E9" , x"ED" , x"ED" , x"E8" , x"CA" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C3" , x"E0" , x"ED" , x"ED" , x"ED" , x"ED" , x"EB" , x"EA" , x"EA" , x"EA" , x"EA" , x"EA" , x"EA" , x"EA" , x"EA" , x"EA" , x"EA" , x"EA" , x"EA" , x"EA" , x"EA" , x"EA" , x"E4" , x"C8" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"C9" , x"E6" , x"ED" , x"ED" , x"ED" , x"ED" , x"EA" , x"C5" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C5" , x"E3" , x"ED" , x"ED" , x"ED" , x"ED" , x"E6" , x"C7" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"CC" , x"E8" , x"ED" , x"ED" , x"ED" , x"C9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C1" , x"E1" , x"ED" , x"ED" , x"ED" , x"D5" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BB" , x"D6" , x"EA" , x"ED" , x"ED" , x"ED" , x"ED" , x"E9" , x"CC" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"C2" , x"D5" , x"E8" , x"EC" , x"ED" , x"ED" , x"ED" , x"EC" , x"EB" , x"EB" , x"EA" , x"EA" , x"EA" , x"EA" , x"EB" , x"EC" , x"ED" , x"ED" , x"ED" , x"ED" , x"E9" , x"D5" , x"BF" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"D4" , x"E9" , x"ED" , x"ED" , x"E8" , x"CA" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"CC" , x"E8" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"E7" , x"CA" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C2" , x"DF" , x"ED" , x"ED" , x"ED" , x"ED" , x"E2" , x"BE" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BA" , x"DA" , x"EC" , x"ED" , x"ED" , x"ED" , x"DF" , x"BE" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"CC" , x"E8" , x"ED" , x"ED" , x"ED" , x"C9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C1" , x"E1" , x"ED" , x"ED" , x"ED" , x"D5" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BE" , x"DD" , x"EB" , x"ED" , x"ED" , x"ED" , x"E9" , x"CC" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BB" , x"CB" , x"DE" , x"E8" , x"EC" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"EC" , x"E9" , x"DF" , x"CA" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"D4" , x"E9" , x"ED" , x"ED" , x"E8" , x"CA" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BA" , x"D3" , x"EB" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"ED" , x"E7" , x"CA" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BC" , x"D8" , x"EB" , x"ED" , x"ED" , x"ED" , x"D8" , x"BA" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"D0" , x"EA" , x"ED" , x"ED" , x"EC" , x"D7" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"CC" , x"E8" , x"ED" , x"ED" , x"ED" , x"C9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C1" , x"E1" , x"ED" , x"ED" , x"ED" , x"D5" , x"BB" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"CA" , x"E4" , x"EC" , x"ED" , x"ED" , x"E9" , x"CC" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B9" , x"C1" , x"CD" , x"DA" , x"E1" , x"E6" , x"E8" , x"EC" , x"EC" , x"ED" , x"ED" , x"ED" , x"EB" , x"E8" , x"E3" , x"DB" , x"CF" , x"C2" , x"BA" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"C6" , x"D2" , x"D4" , x"D4" , x"D1" , x"C0" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BB" , x"C8" , x"D2" , x"D4" , x"D4" , x"D4" , x"D4" , x"D4" , x"D4" , x"D4" , x"D4" , x"D4" , x"D4" , x"D4" , x"D4" , x"D4" , x"D4" , x"D4" , x"D4" , x"D4" , x"D4" , x"D4" , x"D4" , x"CF" , x"C1" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"C5" , x"D3" , x"D4" , x"D4" , x"D4" , x"C4" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C2" , x"D1" , x"D4" , x"D4" , x"D3" , x"C4" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"C2" , x"D1" , x"D4" , x"D4" , x"D4" , x"C1" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BD" , x"CE" , x"D4" , x"D4" , x"D4" , x"C6" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"BC" , x"CB" , x"D3" , x"D4" , x"D4" , x"D2" , x"C3" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"BA" , x"BD" , x"C4" , x"C9" , x"CE" , x"D1" , x"D4" , x"D4" , x"D4" , x"D3" , x"D0" , x"CC" , x"C6" , x"BE" , x"BA" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"B9" , x"B9" , x"B9" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"BA" , x"B9" , x"B9" , x"B9" , x"B9" , x"B9" , x"B9" , x"B9" , x"B9" , x"B9" , x"B9" , x"B9" , x"B9" , x"B9" , x"B9" , x"B9" , x"B9" , x"B9" , x"B9" , x"B9" , x"B9" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"BA" , x"B9" , x"B9" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"B9" , x"B9" , x"B9" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"B9" , x"B9" , x"B9" , x"B9" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"B9" , x"B9" , x"B9" , x"B9" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"BA" , x"B9" , x"B9" , x"B9" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B8" , x"B8" , x"B8" , x"BA" , x"BA" , x"B9" , x"B9" , x"BA" , x"B9" , x"B9" , x"B8" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" ),
( x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" , x"B7" )
);

CONSTANT P2winsG : ImageMatrix(0 TO 99, 0 TO 199) := (
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E4" , x"D3" , x"C8" , x"C0" , x"B7" , x"B7" , x"B7" , x"B8" , x"C1" , x"C7" , x"D2" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"BD" , x"9C" , x"96" , x"96" , x"96" , x"96" , x"96" , x"96" , x"96" , x"96" , x"96" , x"96" , x"96" , x"96" , x"96" , x"96" , x"9A" , x"A5" , x"AE" , x"BC" , x"D5" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E5" , x"C4" , x"9D" , x"96" , x"96" , x"9D" , x"C7" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"CD" , x"9F" , x"96" , x"96" , x"96" , x"96" , x"BF" , x"E5" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DA" , x"A6" , x"97" , x"96" , x"99" , x"B8" , x"E3" , x"E8" , x"E8" , x"E8" , x"C8" , x"9E" , x"96" , x"96" , x"96" , x"CC" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DA" , x"A9" , x"96" , x"96" , x"96" , x"9C" , x"D3" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D2" , x"A4" , x"96" , x"96" , x"9D" , x"C7" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DF" , x"BB" , x"94" , x"6E" , x"54" , x"44" , x"36" , x"34" , x"34" , x"39" , x"46" , x"54" , x"6B" , x"94" , x"B9" , x"D9" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"84" , x"34" , x"29" , x"29" , x"29" , x"29" , x"29" , x"29" , x"29" , x"29" , x"29" , x"29" , x"29" , x"29" , x"29" , x"29" , x"2B" , x"37" , x"3F" , x"4D" , x"68" , x"97" , x"CE" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D9" , x"B2" , x"96" , x"81" , x"78" , x"76" , x"77" , x"8C" , x"A0" , x"BF" , x"DD" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E5" , x"A5" , x"3E" , x"29" , x"29" , x"32" , x"90" , x"E2" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"99" , x"3A" , x"29" , x"29" , x"29" , x"29" , x"6F" , x"D2" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"B6" , x"44" , x"29" , x"29" , x"33" , x"88" , x"DC" , x"E8" , x"E8" , x"E8" , x"9D" , x"3B" , x"29" , x"29" , x"29" , x"A6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C7" , x"55" , x"29" , x"29" , x"29" , x"30" , x"8C" , x"DB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"B2" , x"48" , x"2A" , x"29" , x"38" , x"9B" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E5" , x"C4" , x"83" , x"4C" , x"2E" , x"25" , x"20" , x"1F" , x"1D" , x"1C" , x"1C" , x"1D" , x"1F" , x"20" , x"23" , x"2E" , x"4A" , x"77" , x"BA" , x"E3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"7E" , x"29" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1D" , x"1D" , x"1D" , x"20" , x"2D" , x"4F" , x"9C" , x"DB" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E4" , x"CD" , x"89" , x"52" , x"38" , x"2B" , x"23" , x"20" , x"1F" , x"1F" , x"28" , x"31" , x"3B" , x"64" , x"AE" , x"D8" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"BA" , x"4A" , x"1F" , x"1C" , x"1D" , x"6B" , x"D2" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E4" , x"6A" , x"25" , x"1C" , x"1C" , x"1C" , x"1C" , x"43" , x"B9" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E4" , x"8B" , x"2C" , x"1C" , x"1C" , x"35" , x"A5" , x"E2" , x"E8" , x"E8" , x"E8" , x"99" , x"31" , x"1C" , x"1C" , x"1C" , x"A3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"4A" , x"1C" , x"1C" , x"1C" , x"1D" , x"3E" , x"A5" , x"E0" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"AE" , x"3E" , x"1E" , x"1C" , x"2C" , x"95" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E0" , x"A0" , x"4E" , x"28" , x"1E" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1D" , x"24" , x"45" , x"94" , x"D9" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"7E" , x"29" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1F" , x"34" , x"91" , x"D9" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DF" , x"AE" , x"5F" , x"2D" , x"1F" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"22" , x"3C" , x"80" , x"CB" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CF" , x"66" , x"20" , x"1C" , x"1C" , x"4E" , x"BF" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"47" , x"1E" , x"1C" , x"1C" , x"1C" , x"1C" , x"27" , x"A0" , x"E5" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E2" , x"68" , x"23" , x"1C" , x"1D" , x"4B" , x"C8" , x"E7" , x"E8" , x"E8" , x"E8" , x"99" , x"31" , x"1C" , x"1C" , x"1C" , x"A3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"4A" , x"1C" , x"1C" , x"1C" , x"1C" , x"20" , x"5D" , x"C1" , x"E5" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"AE" , x"3E" , x"1E" , x"1C" , x"2C" , x"95" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E3" , x"A6" , x"44" , x"20" , x"1C" , x"1C" , x"1D" , x"24" , x"34" , x"41" , x"52" , x"56" , x"56" , x"50" , x"43" , x"35" , x"25" , x"1C" , x"1C" , x"1C" , x"1F" , x"37" , x"93" , x"DA" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"7E" , x"29" , x"1C" , x"1C" , x"25" , x"58" , x"73" , x"77" , x"77" , x"77" , x"77" , x"77" , x"77" , x"77" , x"77" , x"77" , x"70" , x"58" , x"43" , x"27" , x"1C" , x"1C" , x"1C" , x"1D" , x"45" , x"AA" , x"E2" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E3" , x"AD" , x"51" , x"25" , x"1D" , x"1C" , x"1C" , x"1F" , x"30" , x"40" , x"44" , x"3A" , x"27" , x"1D" , x"1C" , x"1C" , x"1E" , x"31" , x"77" , x"CD" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E2" , x"84" , x"28" , x"1C" , x"1C" , x"36" , x"B0" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"AB" , x"32" , x"1C" , x"1C" , x"21" , x"1D" , x"1C" , x"1D" , x"78" , x"DB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DA" , x"4B" , x"1F" , x"1C" , x"1F" , x"6E" , x"D5" , x"E8" , x"E8" , x"E8" , x"E8" , x"99" , x"31" , x"1C" , x"1C" , x"1C" , x"A3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"4A" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"2B" , x"82" , x"D8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"AE" , x"3E" , x"1E" , x"1C" , x"2C" , x"95" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C9" , x"5B" , x"21" , x"1C" , x"1C" , x"1E" , x"48" , x"7D" , x"9D" , x"B1" , x"CE" , x"D3" , x"D3" , x"C9" , x"B3" , x"9D" , x"7A" , x"3F" , x"1F" , x"1C" , x"1C" , x"1E" , x"49" , x"AF" , x"E3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"7E" , x"29" , x"1C" , x"1C" , x"2F" , x"9C" , x"D7" , x"DD" , x"DD" , x"DD" , x"DD" , x"DD" , x"DD" , x"DD" , x"DD" , x"DD" , x"DA" , x"C5" , x"B5" , x"86" , x"31" , x"1D" , x"1C" , x"1C" , x"22" , x"65" , x"CB" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"C6" , x"5A" , x"24" , x"1C" , x"1C" , x"20" , x"43" , x"82" , x"A7" , x"B4" , x"B6" , x"AE" , x"98" , x"60" , x"2D" , x"1D" , x"1C" , x"1D" , x"2D" , x"87" , x"DE" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"A2" , x"37" , x"1C" , x"1C" , x"23" , x"9A" , x"E5" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"83" , x"26" , x"1C" , x"1C" , x"4A" , x"29" , x"1C" , x"1C" , x"50" , x"D1" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"BA" , x"37" , x"1C" , x"1C" , x"21" , x"91" , x"DD" , x"E8" , x"E8" , x"E8" , x"E8" , x"99" , x"31" , x"1C" , x"1C" , x"1C" , x"A3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"4A" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1D" , x"3A" , x"AD" , x"E5" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"AE" , x"3E" , x"1E" , x"1C" , x"2C" , x"95" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E3" , x"91" , x"2F" , x"1C" , x"1C" , x"20" , x"5E" , x"B3" , x"DA" , x"E3" , x"E4" , x"E7" , x"E8" , x"E8" , x"E7" , x"E4" , x"E3" , x"D8" , x"AD" , x"4D" , x"21" , x"1C" , x"1C" , x"23" , x"6F" , x"D0" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"7E" , x"29" , x"1C" , x"1C" , x"30" , x"A2" , x"E1" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DF" , x"98" , x"3C" , x"1F" , x"1C" , x"1C" , x"36" , x"9F" , x"E3" , x"E8" , x"E8" , x"E8" , x"E3" , x"7A" , x"29" , x"1C" , x"1C" , x"27" , x"69" , x"BA" , x"E1" , x"E8" , x"E8" , x"E8" , x"E8" , x"E5" , x"D6" , x"9C" , x"42" , x"1E" , x"1C" , x"1C" , x"32" , x"B2" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C2" , x"4C" , x"1C" , x"1C" , x"1C" , x"6F" , x"D9" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D2" , x"5B" , x"1E" , x"1C" , x"31" , x"8A" , x"3D" , x"1D" , x"1C" , x"29" , x"BB" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"92" , x"2A" , x"1C" , x"1C" , x"32" , x"C1" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"99" , x"31" , x"1C" , x"1C" , x"1C" , x"A3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"4A" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1D" , x"51" , x"C7" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"AE" , x"3E" , x"1E" , x"1C" , x"2C" , x"95" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C8" , x"5B" , x"20" , x"1C" , x"1E" , x"50" , x"BD" , x"E5" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"B9" , x"51" , x"21" , x"1C" , x"1C" , x"3B" , x"A8" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"7E" , x"29" , x"1C" , x"1C" , x"30" , x"A2" , x"E1" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D6" , x"7F" , x"29" , x"1C" , x"1C" , x"23" , x"7E" , x"DB" , x"E8" , x"E8" , x"E8" , x"CA" , x"45" , x"1E" , x"1C" , x"1D" , x"5A" , x"BD" , x"E3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DF" , x"97" , x"2F" , x"1C" , x"1C" , x"20" , x"7F" , x"DA" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E3" , x"6B" , x"1F" , x"1C" , x"1C" , x"50" , x"D0" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"B6" , x"43" , x"1C" , x"1C" , x"4B" , x"B5" , x"5B" , x"21" , x"1C" , x"20" , x"8B" , x"DB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E3" , x"70" , x"21" , x"1C" , x"1C" , x"52" , x"D0" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"99" , x"31" , x"1C" , x"1C" , x"1C" , x"A3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"4A" , x"1C" , x"1C" , x"1C" , x"25" , x"1F" , x"1C" , x"1C" , x"26" , x"80" , x"D6" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"AE" , x"3E" , x"1E" , x"1C" , x"2C" , x"95" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"B4" , x"43" , x"1E" , x"1C" , x"28" , x"8A" , x"E0" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DE" , x"8E" , x"31" , x"1D" , x"1C" , x"24" , x"87" , x"DF" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"7E" , x"29" , x"1C" , x"1C" , x"30" , x"A2" , x"E1" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"AF" , x"3E" , x"1E" , x"1C" , x"1D" , x"62" , x"CD" , x"E8" , x"E8" , x"E8" , x"9F" , x"2D" , x"1C" , x"1C" , x"29" , x"A5" , x"E0" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D6" , x"56" , x"20" , x"1C" , x"1D" , x"54" , x"D0" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"8A" , x"27" , x"1C" , x"1C" , x"32" , x"C7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"9A" , x"32" , x"1C" , x"1E" , x"6E" , x"D0" , x"81" , x"29" , x"1C" , x"1F" , x"63" , x"D3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CF" , x"54" , x"1D" , x"1C" , x"1C" , x"7A" , x"DC" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"99" , x"31" , x"1C" , x"1C" , x"1C" , x"A3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"4A" , x"1C" , x"1C" , x"1C" , x"50" , x"34" , x"1E" , x"1C" , x"1D" , x"3E" , x"A6" , x"E2" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"AE" , x"3E" , x"1E" , x"1C" , x"2C" , x"95" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"A7" , x"35" , x"1D" , x"1C" , x"36" , x"A2" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"B8" , x"4D" , x"1F" , x"1C" , x"1D" , x"6A" , x"D4" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"7E" , x"29" , x"1C" , x"1C" , x"30" , x"A2" , x"E1" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C0" , x"52" , x"20" , x"1C" , x"1C" , x"4E" , x"BF" , x"E8" , x"E8" , x"E7" , x"7A" , x"20" , x"1C" , x"1C" , x"48" , x"CB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E4" , x"7F" , x"29" , x"1C" , x"1C" , x"3F" , x"C9" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"B3" , x"34" , x"1C" , x"1C" , x"21" , x"A3" , x"E1" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DB" , x"77" , x"24" , x"1C" , x"29" , x"8E" , x"E0" , x"B2" , x"36" , x"1C" , x"1C" , x"42" , x"BC" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"B1" , x"3F" , x"1C" , x"1C" , x"29" , x"A2" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"99" , x"31" , x"1C" , x"1C" , x"1C" , x"A3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"4A" , x"1C" , x"1C" , x"1C" , x"70" , x"77" , x"2E" , x"1C" , x"1C" , x"21" , x"5A" , x"BF" , x"E5" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"AE" , x"3E" , x"1E" , x"1C" , x"2C" , x"95" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"A4" , x"32" , x"1D" , x"1C" , x"33" , x"9D" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CE" , x"67" , x"33" , x"3F" , x"41" , x"7F" , x"D6" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"7E" , x"29" , x"1C" , x"1C" , x"30" , x"A2" , x"E1" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"56" , x"20" , x"1C" , x"1C" , x"49" , x"BA" , x"E8" , x"E8" , x"DC" , x"6F" , x"2A" , x"26" , x"20" , x"66" , x"D6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"95" , x"2F" , x"1C" , x"1C" , x"37" , x"B1" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DC" , x"4D" , x"1F" , x"1C" , x"1F" , x"7D" , x"D9" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C0" , x"53" , x"1F" , x"1C" , x"3E" , x"AA" , x"E4" , x"CC" , x"54" , x"21" , x"1C" , x"2E" , x"94" , x"DF" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"91" , x"2E" , x"1C" , x"1C" , x"43" , x"BB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"99" , x"31" , x"1C" , x"1C" , x"1C" , x"A3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"4A" , x"1C" , x"1C" , x"1C" , x"77" , x"C0" , x"69" , x"27" , x"1C" , x"1C" , x"26" , x"77" , x"D4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"AE" , x"3E" , x"1E" , x"1C" , x"2C" , x"95" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"AF" , x"3F" , x"1D" , x"1C" , x"21" , x"75" , x"D7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E3" , x"D1" , x"C6" , x"CA" , x"CB" , x"D6" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"7E" , x"29" , x"1C" , x"1C" , x"30" , x"A2" , x"E1" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C0" , x"51" , x"20" , x"1C" , x"1C" , x"54" , x"C2" , x"E8" , x"E8" , x"DC" , x"AC" , x"89" , x"7F" , x"73" , x"9D" , x"DF" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"8D" , x"2C" , x"1C" , x"1C" , x"3B" , x"C0" , x"E5" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E4" , x"6C" , x"25" , x"1C" , x"1E" , x"5C" , x"D2" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"A7" , x"39" , x"1D" , x"1E" , x"58" , x"C8" , x"E6" , x"D7" , x"71" , x"26" , x"1C" , x"24" , x"78" , x"DB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DA" , x"72" , x"23" , x"1C" , x"1C" , x"67" , x"D2" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"99" , x"31" , x"1C" , x"1C" , x"1C" , x"A3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"4A" , x"1C" , x"1C" , x"1C" , x"78" , x"D8" , x"B2" , x"49" , x"1F" , x"1C" , x"1D" , x"35" , x"A1" , x"E2" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"AE" , x"3E" , x"1E" , x"1C" , x"2C" , x"95" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C2" , x"55" , x"1F" , x"1C" , x"1D" , x"39" , x"94" , x"D9" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"7E" , x"29" , x"1C" , x"1C" , x"30" , x"A2" , x"E1" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E5" , x"AC" , x"3C" , x"1E" , x"1C" , x"1C" , x"69" , x"D2" , x"E8" , x"E8" , x"E6" , x"E2" , x"DD" , x"DC" , x"DB" , x"DF" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E4" , x"6A" , x"25" , x"1C" , x"1D" , x"4A" , x"CC" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E5" , x"8E" , x"2C" , x"1C" , x"1C" , x"42" , x"C0" , x"E5" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DC" , x"85" , x"2A" , x"1C" , x"25" , x"79" , x"D9" , x"E8" , x"E3" , x"96" , x"30" , x"1D" , x"1E" , x"58" , x"C7" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C5" , x"57" , x"21" , x"1C" , x"26" , x"8A" , x"E0" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"99" , x"31" , x"1C" , x"1C" , x"1C" , x"A3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"4A" , x"1C" , x"1C" , x"1C" , x"78" , x"DA" , x"DA" , x"8B" , x"30" , x"1C" , x"1C" , x"1F" , x"50" , x"C8" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"AE" , x"3E" , x"1E" , x"1C" , x"2C" , x"95" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DB" , x"7F" , x"28" , x"1C" , x"1C" , x"1F" , x"3B" , x"77" , x"A6" , x"D2" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"7E" , x"29" , x"1C" , x"1C" , x"30" , x"A2" , x"E1" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D3" , x"73" , x"28" , x"1C" , x"1C" , x"26" , x"88" , x"E0" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C0" , x"3D" , x"1E" , x"1C" , x"1E" , x"6D" , x"D5" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"BC" , x"41" , x"1E" , x"1C" , x"32" , x"9F" , x"E1" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D1" , x"5F" , x"23" , x"1C" , x"31" , x"9C" , x"DF" , x"E8" , x"E8" , x"B7" , x"46" , x"1F" , x"1C" , x"3B" , x"A5" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"B4" , x"44" , x"1E" , x"1C" , x"3B" , x"A5" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"99" , x"31" , x"1C" , x"1C" , x"1C" , x"A3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"4A" , x"1C" , x"1C" , x"1C" , x"78" , x"DA" , x"E7" , x"D6" , x"69" , x"22" , x"1C" , x"1C" , x"23" , x"79" , x"D5" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"AE" , x"3E" , x"1E" , x"1C" , x"2C" , x"95" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"C2" , x"54" , x"20" , x"1C" , x"1C" , x"1D" , x"25" , x"35" , x"4E" , x"75" , x"9C" , x"C1" , x"D6" , x"DD" , x"E4" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"7E" , x"29" , x"1C" , x"1C" , x"30" , x"A2" , x"E1" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D4" , x"82" , x"32" , x"1E" , x"1C" , x"1D" , x"44" , x"B0" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DB" , x"78" , x"24" , x"1C" , x"1C" , x"29" , x"A6" , x"E2" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D1" , x"5E" , x"22" , x"1C" , x"27" , x"80" , x"DA" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"BD" , x"43" , x"1F" , x"1C" , x"44" , x"BF" , x"E5" , x"E8" , x"E8" , x"CD" , x"63" , x"20" , x"1C" , x"27" , x"88" , x"DE" , x"E8" , x"E8" , x"E8" , x"E8" , x"E5" , x"9C" , x"2F" , x"1C" , x"1D" , x"54" , x"C0" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"99" , x"31" , x"1C" , x"1C" , x"1C" , x"A3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"4A" , x"1C" , x"1C" , x"1C" , x"78" , x"DA" , x"E8" , x"E8" , x"B8" , x"44" , x"20" , x"1C" , x"1D" , x"37" , x"9A" , x"DD" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"AE" , x"3E" , x"1E" , x"1C" , x"2C" , x"95" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E4" , x"AE" , x"4D" , x"22" , x"1C" , x"1C" , x"1C" , x"1C" , x"1D" , x"25" , x"2E" , x"3D" , x"52" , x"70" , x"95" , x"B7" , x"C8" , x"DA" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"7E" , x"29" , x"1C" , x"1C" , x"30" , x"A2" , x"E1" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"CF" , x"BD" , x"A6" , x"74" , x"32" , x"1E" , x"1C" , x"1C" , x"26" , x"79" , x"D6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DD" , x"98" , x"3B" , x"1D" , x"1C" , x"1D" , x"5C" , x"D0" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DA" , x"7B" , x"27" , x"1C" , x"20" , x"66" , x"D2" , x"E7" , x"E8" , x"E8" , x"E8" , x"E5" , x"96" , x"30" , x"1C" , x"1F" , x"67" , x"D1" , x"E8" , x"E8" , x"E8" , x"E1" , x"82" , x"27" , x"1C" , x"1E" , x"64" , x"CE" , x"E8" , x"E8" , x"E8" , x"E8" , x"D9" , x"78" , x"27" , x"1C" , x"22" , x"73" , x"D7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"99" , x"31" , x"1C" , x"1C" , x"1C" , x"A3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"4A" , x"1C" , x"1C" , x"1C" , x"78" , x"DA" , x"E8" , x"E8" , x"DF" , x"90" , x"34" , x"1E" , x"1C" , x"21" , x"53" , x"BA" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"AE" , x"3E" , x"1E" , x"1C" , x"2C" , x"95" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E0" , x"AE" , x"61" , x"2C" , x"1D" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1D" , x"20" , x"26" , x"2E" , x"3E" , x"59" , x"79" , x"A2" , x"C6" , x"E1" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"7E" , x"29" , x"1C" , x"1C" , x"25" , x"56" , x"70" , x"74" , x"74" , x"74" , x"74" , x"74" , x"74" , x"74" , x"74" , x"74" , x"5D" , x"4C" , x"39" , x"27" , x"1D" , x"1C" , x"1C" , x"1D" , x"4D" , x"B9" , x"E3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E3" , x"A9" , x"4B" , x"21" , x"1C" , x"1C" , x"37" , x"A0" , x"E3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E3" , x"9F" , x"34" , x"1D" , x"1C" , x"4C" , x"BD" , x"E5" , x"E8" , x"E8" , x"E8" , x"E4" , x"70" , x"26" , x"1C" , x"20" , x"8D" , x"DC" , x"E8" , x"E8" , x"E8" , x"E7" , x"A2" , x"37" , x"1C" , x"1C" , x"43" , x"BB" , x"E8" , x"E8" , x"E8" , x"E8" , x"CE" , x"5A" , x"21" , x"1C" , x"2C" , x"8F" , x"DE" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"99" , x"31" , x"1C" , x"1C" , x"1C" , x"A3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"4A" , x"1C" , x"1C" , x"1C" , x"78" , x"DA" , x"E8" , x"E8" , x"E8" , x"CD" , x"68" , x"24" , x"1C" , x"1C" , x"28" , x"78" , x"D4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"AE" , x"3E" , x"1E" , x"1C" , x"2C" , x"95" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E2" , x"C5" , x"93" , x"51" , x"26" , x"1D" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1E" , x"20" , x"26" , x"37" , x"56" , x"8A" , x"CA" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"7E" , x"29" , x"1C" , x"1C" , x"1C" , x"1D" , x"1E" , x"1E" , x"1E" , x"1E" , x"1E" , x"1E" , x"1E" , x"1E" , x"1E" , x"1E" , x"1D" , x"1D" , x"1C" , x"1C" , x"1C" , x"1C" , x"21" , x"4D" , x"B8" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E2" , x"A2" , x"47" , x"21" , x"1C" , x"1D" , x"34" , x"8E" , x"DA" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"BD" , x"4F" , x"1F" , x"1C" , x"37" , x"A1" , x"E4" , x"E8" , x"E8" , x"E8" , x"D1" , x"43" , x"1E" , x"1C" , x"2B" , x"BC" , x"E5" , x"E8" , x"E8" , x"E8" , x"E8" , x"C5" , x"4D" , x"1C" , x"1C" , x"26" , x"A1" , x"E6" , x"E8" , x"E8" , x"E7" , x"BD" , x"3C" , x"1D" , x"1C" , x"3E" , x"B9" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"99" , x"31" , x"1C" , x"1C" , x"1C" , x"A3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"4A" , x"1C" , x"1C" , x"1C" , x"78" , x"DA" , x"E8" , x"E8" , x"E8" , x"E4" , x"B6" , x"50" , x"21" , x"1C" , x"1C" , x"2D" , x"9A" , x"E2" , x"E8" , x"E8" , x"E8" , x"E8" , x"AE" , x"3E" , x"1E" , x"1C" , x"2C" , x"95" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"E2" , x"CF" , x"B2" , x"7E" , x"52" , x"35" , x"29" , x"22" , x"1D" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1E" , x"29" , x"4D" , x"9E" , x"D8" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"7E" , x"29" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"21" , x"37" , x"65" , x"B4" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DB" , x"A4" , x"43" , x"20" , x"1C" , x"1C" , x"2F" , x"7A" , x"CC" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D0" , x"66" , x"20" , x"1C" , x"29" , x"8D" , x"E2" , x"E8" , x"E8" , x"E8" , x"AA" , x"32" , x"1C" , x"1C" , x"4D" , x"CF" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E3" , x"6D" , x"20" , x"1C" , x"1D" , x"73" , x"DA" , x"E8" , x"E8" , x"E4" , x"93" , x"2D" , x"1C" , x"1E" , x"5B" , x"D1" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"99" , x"31" , x"1C" , x"1C" , x"1C" , x"A3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"4A" , x"1C" , x"1C" , x"1C" , x"78" , x"DA" , x"E8" , x"E8" , x"E8" , x"E8" , x"E2" , x"99" , x"33" , x"1C" , x"1C" , x"1D" , x"4A" , x"BE" , x"E4" , x"E8" , x"E8" , x"E8" , x"AE" , x"3E" , x"1E" , x"1C" , x"2C" , x"95" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E5" , x"DA" , x"CF" , x"B1" , x"8E" , x"70" , x"54" , x"3D" , x"2B" , x"20" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1F" , x"3C" , x"8F" , x"D5" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"7E" , x"29" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"26" , x"32" , x"3F" , x"55" , x"7A" , x"A3" , x"C9" , x"E3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D9" , x"93" , x"44" , x"1F" , x"1C" , x"1C" , x"28" , x"7A" , x"CA" , x"E3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E2" , x"87" , x"29" , x"1C" , x"1E" , x"70" , x"D6" , x"E8" , x"E8" , x"E8" , x"84" , x"26" , x"1C" , x"1C" , x"76" , x"DB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"92" , x"2A" , x"1C" , x"1C" , x"4C" , x"CF" , x"E8" , x"E8" , x"E4" , x"6F" , x"26" , x"1C" , x"20" , x"81" , x"DA" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"99" , x"31" , x"1C" , x"1C" , x"1C" , x"A3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"4A" , x"1C" , x"1C" , x"1C" , x"78" , x"DA" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D2" , x"6B" , x"23" , x"1C" , x"1C" , x"24" , x"74" , x"D2" , x"E7" , x"E8" , x"E8" , x"AE" , x"3E" , x"1E" , x"1C" , x"2C" , x"95" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E3" , x"DE" , x"D8" , x"C7" , x"AB" , x"90" , x"73" , x"50" , x"2E" , x"1D" , x"1C" , x"1C" , x"1C" , x"1F" , x"3E" , x"A1" , x"E2" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"7E" , x"29" , x"1C" , x"1C" , x"29" , x"6F" , x"95" , x"9B" , x"9B" , x"9B" , x"9B" , x"9B" , x"9B" , x"9B" , x"9B" , x"9B" , x"A0" , x"AB" , x"B4" , x"C4" , x"DA" , x"E4" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D7" , x"85" , x"3B" , x"20" , x"1C" , x"1D" , x"28" , x"72" , x"CE" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"A6" , x"3B" , x"1C" , x"1C" , x"4F" , x"C1" , x"E8" , x"E8" , x"DB" , x"63" , x"1F" , x"1C" , x"27" , x"9E" , x"E5" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"B9" , x"36" , x"1C" , x"1C" , x"2B" , x"BA" , x"E6" , x"E8" , x"DF" , x"4D" , x"1F" , x"1C" , x"27" , x"B1" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"99" , x"31" , x"1C" , x"1C" , x"1C" , x"A3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"4A" , x"1C" , x"1C" , x"1C" , x"78" , x"DA" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"C1" , x"45" , x"1F" , x"1C" , x"1D" , x"37" , x"9A" , x"DF" , x"E8" , x"E8" , x"AE" , x"3E" , x"1E" , x"1C" , x"2C" , x"95" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"E4" , x"E1" , x"D7" , x"C0" , x"A4" , x"61" , x"2D" , x"1F" , x"1C" , x"1C" , x"20" , x"58" , x"C9" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"7E" , x"29" , x"1C" , x"1C" , x"30" , x"A2" , x"E1" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E3" , x"C4" , x"61" , x"2B" , x"1E" , x"1C" , x"1E" , x"3B" , x"8F" , x"D4" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C8" , x"50" , x"1C" , x"1C" , x"36" , x"B0" , x"E8" , x"E8" , x"B7" , x"43" , x"1C" , x"1C" , x"42" , x"B9" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DD" , x"52" , x"20" , x"1C" , x"20" , x"91" , x"DC" , x"E8" , x"B8" , x"36" , x"1C" , x"1C" , x"45" , x"CC" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"99" , x"31" , x"1C" , x"1C" , x"1C" , x"A3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"4A" , x"1C" , x"1C" , x"1C" , x"78" , x"DA" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E4" , x"97" , x"37" , x"1E" , x"1C" , x"1F" , x"4A" , x"B2" , x"E3" , x"E8" , x"AE" , x"3E" , x"1E" , x"1C" , x"2C" , x"95" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"D1" , x"9A" , x"46" , x"20" , x"1C" , x"1C" , x"25" , x"9C" , x"E3" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"7E" , x"29" , x"1C" , x"1C" , x"30" , x"A2" , x"E1" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DD" , x"AC" , x"59" , x"25" , x"1D" , x"1C" , x"1D" , x"44" , x"94" , x"D6" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E4" , x"6E" , x"21" , x"1C" , x"22" , x"97" , x"E3" , x"E8" , x"9B" , x"32" , x"1C" , x"1D" , x"66" , x"CF" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E4" , x"77" , x"29" , x"1C" , x"1F" , x"72" , x"D6" , x"E8" , x"99" , x"2C" , x"1C" , x"1C" , x"69" , x"D6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"99" , x"31" , x"1C" , x"1C" , x"1C" , x"A3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"4A" , x"1C" , x"1C" , x"1C" , x"78" , x"DA" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"D1" , x"75" , x"2A" , x"1C" , x"1C" , x"24" , x"6C" , x"D1" , x"E8" , x"AE" , x"3E" , x"1E" , x"1C" , x"2C" , x"95" , x"E4" , x"E8" , x"E8" , x"E8" , x"E6" , x"D0" , x"B9" , x"B2" , x"AD" , x"B8" , x"E0" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"DA" , x"8E" , x"31" , x"1C" , x"1C" , x"1D" , x"74" , x"D9" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"7E" , x"29" , x"1C" , x"1C" , x"30" , x"A2" , x"E1" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DD" , x"9A" , x"4B" , x"24" , x"1C" , x"1C" , x"1E" , x"48" , x"A7" , x"DA" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"91" , x"29" , x"1C" , x"1C" , x"73" , x"DB" , x"DC" , x"7A" , x"24" , x"1C" , x"27" , x"89" , x"DF" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E5" , x"9C" , x"30" , x"1C" , x"1E" , x"52" , x"D0" , x"E8" , x"7A" , x"22" , x"1C" , x"21" , x"94" , x"E3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"99" , x"31" , x"1C" , x"1C" , x"1C" , x"A3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"4A" , x"1C" , x"1C" , x"1C" , x"78" , x"DA" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"B9" , x"50" , x"1F" , x"1C" , x"1C" , x"30" , x"97" , x"E1" , x"AE" , x"3E" , x"1E" , x"1C" , x"2C" , x"95" , x"E4" , x"E8" , x"E8" , x"E8" , x"E3" , x"91" , x"4E" , x"40" , x"39" , x"5A" , x"CA" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"CC" , x"4C" , x"1C" , x"1C" , x"1C" , x"5F" , x"D3" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"7E" , x"29" , x"1C" , x"1C" , x"30" , x"A2" , x"E1" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"E0" , x"8B" , x"3C" , x"21" , x"1C" , x"1D" , x"28" , x"5B" , x"AE" , x"E0" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"B6" , x"35" , x"1C" , x"1C" , x"53" , x"D1" , x"C6" , x"5A" , x"21" , x"1C" , x"39" , x"A3" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C1" , x"48" , x"20" , x"1C" , x"3A" , x"B2" , x"CE" , x"59" , x"1D" , x"1C" , x"36" , x"B1" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"99" , x"31" , x"1C" , x"1C" , x"1C" , x"A3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"4A" , x"1C" , x"1C" , x"1C" , x"78" , x"DA" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E0" , x"99" , x"37" , x"1D" , x"1C" , x"1D" , x"43" , x"BD" , x"AB" , x"3E" , x"1E" , x"1C" , x"2C" , x"95" , x"E4" , x"E8" , x"E8" , x"E8" , x"E2" , x"82" , x"2B" , x"1E" , x"1D" , x"3A" , x"AB" , x"E3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"67" , x"20" , x"1C" , x"1C" , x"53" , x"D0" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"7E" , x"29" , x"1C" , x"1C" , x"30" , x"A2" , x"E1" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"CD" , x"7D" , x"30" , x"1D" , x"1C" , x"1C" , x"34" , x"7B" , x"C3" , x"E3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DC" , x"4E" , x"1F" , x"1C" , x"36" , x"C4" , x"B2" , x"40" , x"1E" , x"1D" , x"53" , x"C3" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"6C" , x"25" , x"1C" , x"2E" , x"94" , x"AB" , x"42" , x"1C" , x"1C" , x"59" , x"C8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"99" , x"31" , x"1C" , x"1C" , x"1C" , x"A3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"4A" , x"1C" , x"1C" , x"1C" , x"78" , x"DA" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DD" , x"79" , x"25" , x"1C" , x"1C" , x"20" , x"6A" , x"94" , x"3C" , x"1E" , x"1C" , x"2C" , x"95" , x"E4" , x"E8" , x"E8" , x"E8" , x"E5" , x"9E" , x"31" , x"1C" , x"1C" , x"29" , x"82" , x"D9" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E4" , x"63" , x"20" , x"1C" , x"1C" , x"5F" , x"D3" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"7E" , x"29" , x"1C" , x"1C" , x"30" , x"A2" , x"E1" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D2" , x"7A" , x"32" , x"1D" , x"1C" , x"1C" , x"37" , x"8C" , x"D0" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E3" , x"72" , x"26" , x"1C" , x"24" , x"A5" , x"93" , x"2E" , x"1C" , x"23" , x"73" , x"D7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E1" , x"8E" , x"2C" , x"1C" , x"28" , x"81" , x"8F" , x"32" , x"1C" , x"20" , x"7A" , x"DA" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"99" , x"31" , x"1C" , x"1C" , x"1C" , x"A3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"4A" , x"1C" , x"1C" , x"1C" , x"78" , x"DA" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"BF" , x"4C" , x"20" , x"1C" , x"1C" , x"32" , x"59" , x"33" , x"1D" , x"1C" , x"2C" , x"95" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"C0" , x"44" , x"1E" , x"1C" , x"1E" , x"4D" , x"B9" , x"E5" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C6" , x"4A" , x"1C" , x"1C" , x"1C" , x"71" , x"D9" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"7E" , x"29" , x"1C" , x"1C" , x"30" , x"A2" , x"E1" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DB" , x"89" , x"36" , x"1F" , x"1C" , x"1E" , x"43" , x"96" , x"D9" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E5" , x"97" , x"2E" , x"1C" , x"21" , x"77" , x"68" , x"27" , x"1C" , x"2D" , x"93" , x"DE" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"AE" , x"3E" , x"1D" , x"21" , x"65" , x"71" , x"27" , x"1C" , x"30" , x"99" , x"E3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"99" , x"31" , x"1C" , x"1C" , x"1C" , x"A3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"4A" , x"1C" , x"1C" , x"1C" , x"78" , x"DA" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E3" , x"9C" , x"38" , x"1E" , x"1C" , x"20" , x"29" , x"24" , x"1C" , x"1C" , x"2C" , x"95" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"71" , x"24" , x"1C" , x"1C" , x"29" , x"6C" , x"CE" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DC" , x"8B" , x"2F" , x"1C" , x"1C" , x"25" , x"9B" , x"E2" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"7E" , x"29" , x"1C" , x"1C" , x"30" , x"A2" , x"E1" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E3" , x"95" , x"39" , x"1F" , x"1C" , x"21" , x"4B" , x"A7" , x"DC" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C0" , x"42" , x"1E" , x"1F" , x"51" , x"41" , x"20" , x"1C" , x"3D" , x"B8" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C6" , x"5A" , x"21" , x"1C" , x"3F" , x"48" , x"20" , x"1C" , x"48" , x"B6" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"99" , x"31" , x"1C" , x"1C" , x"1C" , x"A3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"4A" , x"1C" , x"1C" , x"1C" , x"78" , x"DA" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"78" , x"29" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"2C" , x"95" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E4" , x"AD" , x"43" , x"1F" , x"1C" , x"1C" , x"27" , x"64" , x"BC" , x"DC" , x"E5" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E5" , x"D3" , x"8F" , x"3C" , x"1F" , x"1C" , x"1E" , x"51" , x"C4" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"7E" , x"29" , x"1C" , x"1C" , x"30" , x"A2" , x"E1" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C0" , x"47" , x"1F" , x"1C" , x"1C" , x"40" , x"A3" , x"DC" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D0" , x"5F" , x"22" , x"1D" , x"2F" , x"24" , x"1D" , x"1E" , x"60" , x"D1" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DB" , x"79" , x"25" , x"1C" , x"29" , x"2D" , x"1E" , x"21" , x"68" , x"D3" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"99" , x"31" , x"1C" , x"1C" , x"1C" , x"A3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"4A" , x"1C" , x"1C" , x"1C" , x"78" , x"DA" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E5" , x"C0" , x"5B" , x"21" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"2C" , x"95" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DA" , x"87" , x"2E" , x"1C" , x"1C" , x"1C" , x"24" , x"44" , x"7D" , x"AE" , x"C8" , x"D5" , x"E3" , x"E7" , x"E7" , x"E0" , x"D3" , x"C7" , x"AA" , x"6B" , x"32" , x"1E" , x"1C" , x"1D" , x"37" , x"9A" , x"E0" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"7E" , x"29" , x"1C" , x"1C" , x"30" , x"A2" , x"E1" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DF" , x"81" , x"27" , x"1C" , x"1C" , x"1C" , x"48" , x"82" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"9C" , x"CC" , x"E6" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DB" , x"82" , x"28" , x"1C" , x"1F" , x"1D" , x"1C" , x"1F" , x"87" , x"DA" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"9A" , x"33" , x"1C" , x"1E" , x"1E" , x"1C" , x"29" , x"84" , x"DB" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"99" , x"31" , x"1C" , x"1C" , x"1C" , x"A3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"4A" , x"1C" , x"1C" , x"1C" , x"78" , x"DA" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E3" , x"A2" , x"39" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"2C" , x"95" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"CE" , x"6B" , x"27" , x"1D" , x"1C" , x"1C" , x"1F" , x"29" , x"3E" , x"59" , x"72" , x"89" , x"91" , x"91" , x"84" , x"6C" , x"56" , x"39" , x"25" , x"1E" , x"1C" , x"1D" , x"2D" , x"7B" , x"CE" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"7E" , x"29" , x"1C" , x"1C" , x"30" , x"A2" , x"E1" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"BB" , x"4D" , x"1D" , x"1C" , x"1C" , x"1C" , x"20" , x"27" , x"27" , x"27" , x"27" , x"27" , x"27" , x"27" , x"27" , x"27" , x"27" , x"27" , x"27" , x"27" , x"27" , x"27" , x"3D" , x"A9" , x"E2" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E5" , x"A4" , x"34" , x"1D" , x"1C" , x"1C" , x"1C" , x"24" , x"B1" , x"E3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"B9" , x"44" , x"1C" , x"1C" , x"1C" , x"1C" , x"34" , x"A5" , x"E2" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"99" , x"31" , x"1C" , x"1C" , x"1C" , x"A3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"4A" , x"1C" , x"1C" , x"1C" , x"78" , x"DA" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D9" , x"75" , x"25" , x"1C" , x"1C" , x"1C" , x"1C" , x"2C" , x"95" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"C3" , x"70" , x"2D" , x"1E" , x"1C" , x"1C" , x"1C" , x"1E" , x"20" , x"24" , x"27" , x"27" , x"27" , x"26" , x"23" , x"20" , x"1D" , x"1C" , x"1C" , x"1C" , x"29" , x"79" , x"C9" , x"E3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"7E" , x"29" , x"1C" , x"1C" , x"30" , x"A2" , x"E1" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"95" , x"2E" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"32" , x"A5" , x"E2" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"BE" , x"4E" , x"20" , x"1C" , x"1C" , x"1C" , x"47" , x"CD" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E1" , x"63" , x"1E" , x"1C" , x"1C" , x"1D" , x"4E" , x"CA" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"99" , x"31" , x"1C" , x"1C" , x"1C" , x"A3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"4A" , x"1C" , x"1C" , x"1C" , x"78" , x"DA" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D0" , x"56" , x"21" , x"1C" , x"1C" , x"1C" , x"2C" , x"95" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"D4" , x"9C" , x"54" , x"2D" , x"20" , x"1D" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"20" , x"2A" , x"4F" , x"9D" , x"D7" , x"E5" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"7E" , x"29" , x"1C" , x"1C" , x"30" , x"A2" , x"E1" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DC" , x"7B" , x"25" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"1C" , x"32" , x"A5" , x"E2" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"6E" , x"21" , x"1C" , x"1C" , x"1C" , x"6F" , x"D9" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"87" , x"28" , x"1C" , x"1C" , x"20" , x"72" , x"D7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"99" , x"31" , x"1C" , x"1C" , x"1C" , x"A3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"C4" , x"4A" , x"1C" , x"1C" , x"1C" , x"78" , x"DA" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E5" , x"A0" , x"3D" , x"1E" , x"1C" , x"1C" , x"2C" , x"95" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"DF" , x"C4" , x"95" , x"67" , x"48" , x"3A" , x"2D" , x"25" , x"1E" , x"1C" , x"1C" , x"1F" , x"26" , x"30" , x"42" , x"64" , x"91" , x"C0" , x"DF" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"AF" , x"82" , x"7A" , x"7A" , x"85" , x"C2" , x"E3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"DD" , x"A6" , x"7F" , x"7A" , x"7A" , x"7A" , x"7A" , x"7A" , x"7A" , x"7A" , x"7A" , x"7A" , x"7A" , x"7A" , x"7A" , x"7A" , x"7A" , x"7A" , x"7A" , x"7A" , x"7A" , x"7A" , x"7A" , x"86" , x"C4" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E5" , x"B1" , x"80" , x"7A" , x"7A" , x"7A" , x"B5" , x"E3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"BF" , x"84" , x"7A" , x"7A" , x"7D" , x"B4" , x"E1" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"BE" , x"87" , x"7A" , x"7A" , x"7A" , x"C3" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D5" , x"94" , x"7A" , x"7A" , x"7A" , x"AC" , x"E1" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"D7" , x"9C" , x"7E" , x"7A" , x"7A" , x"83" , x"BC" , x"E5" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E5" , x"DF" , x"D2" , x"B8" , x"A5" , x"94" , x"87" , x"7D" , x"7A" , x"7A" , x"7E" , x"89" , x"98" , x"B0" , x"D3" , x"DE" , x"E5" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E4" , x"E0" , x"DF" , x"DF" , x"E0" , x"E5" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"E3" , x"E0" , x"DF" , x"DF" , x"DF" , x"DF" , x"DF" , x"DF" , x"DF" , x"DF" , x"DF" , x"DF" , x"DF" , x"DF" , x"DF" , x"DF" , x"DF" , x"DF" , x"DF" , x"DF" , x"DF" , x"DF" , x"E0" , x"E5" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E4" , x"E0" , x"DF" , x"DF" , x"DF" , x"E4" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E5" , x"E0" , x"DF" , x"DF" , x"DF" , x"E4" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E5" , x"E0" , x"DF" , x"DF" , x"DF" , x"E5" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E6" , x"E2" , x"DF" , x"DF" , x"DF" , x"E4" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"E3" , x"E0" , x"DF" , x"DF" , x"E0" , x"E5" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E7" , x"E5" , x"E4" , x"E2" , x"E1" , x"E0" , x"DF" , x"DF" , x"E0" , x"E1" , x"E3" , x"E5" , x"E7" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" ),
( x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" , x"E8" )
);

CONSTANT P2winsB : ImageMatrix(0 TO 99, 0 TO 199) := (
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"90" , x"87" , x"81" , x"7C" , x"78" , x"78" , x"78" , x"78" , x"7C" , x"80" , x"87" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"7A" , x"68" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"68" , x"6E" , x"72" , x"7B" , x"87" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"7E" , x"69" , x"66" , x"66" , x"6A" , x"80" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"83" , x"6B" , x"66" , x"66" , x"66" , x"66" , x"7B" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8B" , x"6F" , x"66" , x"66" , x"67" , x"79" , x"8F" , x"92" , x"92" , x"92" , x"81" , x"6A" , x"66" , x"66" , x"66" , x"83" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8B" , x"70" , x"66" , x"66" , x"66" , x"69" , x"87" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"86" , x"6D" , x"66" , x"66" , x"69" , x"81" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8E" , x"7A" , x"64" , x"4F" , x"42" , x"39" , x"32" , x"31" , x"31" , x"34" , x"3A" , x"42" , x"4F" , x"65" , x"79" , x"8A" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"5B" , x"32" , x"2B" , x"2B" , x"2B" , x"2B" , x"2B" , x"2B" , x"2B" , x"2B" , x"2B" , x"2B" , x"2B" , x"2B" , x"2B" , x"2B" , x"2C" , x"32" , x"36" , x"3F" , x"4C" , x"66" , x"83" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"89" , x"75" , x"66" , x"5B" , x"55" , x"54" , x"55" , x"60" , x"6B" , x"7B" , x"8C" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"90" , x"6D" , x"36" , x"2C" , x"2B" , x"2F" , x"62" , x"8E" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"68" , x"34" , x"2B" , x"2B" , x"2B" , x"2B" , x"51" , x"86" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"77" , x"3A" , x"2C" , x"2B" , x"31" , x"5E" , x"8B" , x"92" , x"92" , x"92" , x"6A" , x"35" , x"2B" , x"2B" , x"2B" , x"6F" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"80" , x"43" , x"2B" , x"2B" , x"2B" , x"2E" , x"62" , x"8B" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"75" , x"3C" , x"2C" , x"2B" , x"33" , x"68" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"7F" , x"5C" , x"3F" , x"2D" , x"28" , x"26" , x"25" , x"25" , x"24" , x"24" , x"25" , x"25" , x"26" , x"28" , x"2D" , x"3D" , x"55" , x"79" , x"8F" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"58" , x"2B" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"25" , x"25" , x"25" , x"26" , x"2D" , x"40" , x"6A" , x"8B" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"90" , x"84" , x"5D" , x"42" , x"33" , x"2D" , x"28" , x"26" , x"26" , x"26" , x"2A" , x"2F" , x"34" , x"4B" , x"72" , x"8A" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7A" , x"3D" , x"26" , x"24" , x"25" , x"4F" , x"86" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"90" , x"4F" , x"28" , x"24" , x"24" , x"24" , x"24" , x"39" , x"79" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"60" , x"2C" , x"24" , x"24" , x"32" , x"6E" , x"8E" , x"92" , x"92" , x"92" , x"67" , x"2F" , x"24" , x"24" , x"24" , x"6D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7F" , x"3D" , x"24" , x"24" , x"24" , x"25" , x"37" , x"6E" , x"8D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"73" , x"37" , x"25" , x"24" , x"2C" , x"65" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8E" , x"6B" , x"40" , x"2B" , x"25" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"25" , x"29" , x"3A" , x"65" , x"89" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"58" , x"2B" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"25" , x"31" , x"63" , x"8A" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8E" , x"72" , x"48" , x"2D" , x"25" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"28" , x"36" , x"5A" , x"82" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"84" , x"4B" , x"26" , x"24" , x"24" , x"40" , x"7C" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"87" , x"3C" , x"25" , x"24" , x"24" , x"24" , x"24" , x"2A" , x"6A" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8E" , x"4D" , x"28" , x"24" , x"25" , x"3E" , x"80" , x"91" , x"92" , x"92" , x"92" , x"67" , x"2F" , x"24" , x"24" , x"24" , x"6D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7F" , x"3D" , x"24" , x"24" , x"24" , x"24" , x"26" , x"47" , x"7E" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"73" , x"37" , x"25" , x"24" , x"2C" , x"65" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8F" , x"6F" , x"39" , x"26" , x"24" , x"24" , x"25" , x"28" , x"31" , x"38" , x"41" , x"44" , x"44" , x"3F" , x"38" , x"31" , x"28" , x"24" , x"24" , x"24" , x"25" , x"32" , x"65" , x"8B" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"58" , x"2B" , x"24" , x"24" , x"28" , x"44" , x"53" , x"55" , x"55" , x"55" , x"55" , x"55" , x"55" , x"55" , x"55" , x"55" , x"52" , x"44" , x"38" , x"29" , x"24" , x"24" , x"24" , x"25" , x"3A" , x"70" , x"8E" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8F" , x"73" , x"41" , x"29" , x"25" , x"24" , x"24" , x"25" , x"2E" , x"37" , x"39" , x"34" , x"2A" , x"24" , x"24" , x"24" , x"25" , x"2F" , x"55" , x"84" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8E" , x"5D" , x"2B" , x"24" , x"24" , x"33" , x"74" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"71" , x"30" , x"24" , x"24" , x"27" , x"24" , x"24" , x"25" , x"56" , x"8B" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8A" , x"3D" , x"26" , x"24" , x"25" , x"4F" , x"88" , x"92" , x"92" , x"92" , x"92" , x"67" , x"2F" , x"24" , x"24" , x"24" , x"6D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7F" , x"3D" , x"24" , x"24" , x"24" , x"24" , x"24" , x"2C" , x"5C" , x"8A" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"73" , x"37" , x"25" , x"24" , x"2C" , x"65" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"80" , x"46" , x"26" , x"24" , x"24" , x"25" , x"3B" , x"58" , x"6A" , x"74" , x"84" , x"87" , x"87" , x"81" , x"75" , x"6A" , x"58" , x"36" , x"25" , x"24" , x"24" , x"25" , x"3C" , x"73" , x"8F" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"58" , x"2B" , x"24" , x"24" , x"2E" , x"69" , x"89" , x"8D" , x"8D" , x"8D" , x"8D" , x"8D" , x"8D" , x"8D" , x"8D" , x"8D" , x"8A" , x"7F" , x"76" , x"5E" , x"30" , x"25" , x"24" , x"24" , x"27" , x"4C" , x"83" , x"91" , x"92" , x"92" , x"92" , x"92" , x"7F" , x"46" , x"28" , x"24" , x"24" , x"26" , x"38" , x"5B" , x"6F" , x"77" , x"77" , x"73" , x"67" , x"49" , x"2E" , x"25" , x"24" , x"25" , x"2D" , x"5F" , x"8D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"6C" , x"32" , x"24" , x"24" , x"28" , x"67" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"5B" , x"29" , x"24" , x"24" , x"3C" , x"2B" , x"24" , x"24" , x"40" , x"86" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"79" , x"32" , x"24" , x"24" , x"27" , x"63" , x"8D" , x"92" , x"92" , x"92" , x"92" , x"67" , x"2F" , x"24" , x"24" , x"24" , x"6D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7F" , x"3D" , x"24" , x"24" , x"24" , x"24" , x"24" , x"25" , x"34" , x"72" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"73" , x"37" , x"25" , x"24" , x"2C" , x"65" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8F" , x"62" , x"2F" , x"24" , x"24" , x"26" , x"48" , x"75" , x"8B" , x"8F" , x"90" , x"91" , x"92" , x"92" , x"91" , x"91" , x"8F" , x"8A" , x"72" , x"3F" , x"27" , x"24" , x"24" , x"28" , x"51" , x"85" , x"91" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"58" , x"2B" , x"24" , x"24" , x"2E" , x"6C" , x"8E" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8D" , x"67" , x"35" , x"26" , x"24" , x"24" , x"33" , x"6B" , x"8F" , x"92" , x"92" , x"92" , x"8F" , x"57" , x"2B" , x"24" , x"24" , x"29" , x"4E" , x"79" , x"8E" , x"92" , x"92" , x"92" , x"92" , x"90" , x"88" , x"69" , x"38" , x"25" , x"24" , x"24" , x"2F" , x"76" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7E" , x"3E" , x"24" , x"24" , x"24" , x"50" , x"89" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"87" , x"46" , x"25" , x"24" , x"2F" , x"5E" , x"36" , x"25" , x"24" , x"2B" , x"7A" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"63" , x"2B" , x"24" , x"24" , x"31" , x"7C" , x"92" , x"92" , x"92" , x"92" , x"92" , x"67" , x"2F" , x"24" , x"24" , x"24" , x"6D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7F" , x"3D" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"25" , x"41" , x"80" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"73" , x"37" , x"25" , x"24" , x"2C" , x"65" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"81" , x"46" , x"26" , x"24" , x"25" , x"40" , x"7A" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"78" , x"40" , x"26" , x"24" , x"24" , x"35" , x"6F" , x"91" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"58" , x"2B" , x"24" , x"24" , x"2E" , x"6C" , x"8E" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"88" , x"59" , x"2C" , x"24" , x"24" , x"28" , x"58" , x"8A" , x"92" , x"92" , x"92" , x"82" , x"3A" , x"25" , x"24" , x"25" , x"46" , x"7B" , x"8F" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8E" , x"66" , x"2E" , x"24" , x"24" , x"26" , x"59" , x"8A" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8F" , x"4F" , x"25" , x"24" , x"24" , x"40" , x"85" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"78" , x"3A" , x"24" , x"24" , x"3D" , x"76" , x"46" , x"27" , x"24" , x"26" , x"60" , x"8B" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8F" , x"52" , x"27" , x"24" , x"24" , x"41" , x"85" , x"92" , x"92" , x"92" , x"92" , x"92" , x"67" , x"2F" , x"24" , x"24" , x"24" , x"6D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7F" , x"3D" , x"24" , x"24" , x"24" , x"29" , x"26" , x"24" , x"24" , x"29" , x"5A" , x"89" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"73" , x"37" , x"25" , x"24" , x"2C" , x"65" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"76" , x"3A" , x"25" , x"24" , x"2B" , x"60" , x"8E" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8D" , x"62" , x"2F" , x"25" , x"24" , x"29" , x"5E" , x"8D" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"58" , x"2B" , x"24" , x"24" , x"2E" , x"6C" , x"8E" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"73" , x"37" , x"25" , x"24" , x"25" , x"4A" , x"84" , x"92" , x"92" , x"92" , x"6B" , x"2E" , x"24" , x"24" , x"2B" , x"6E" , x"8E" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"88" , x"42" , x"26" , x"24" , x"25" , x"42" , x"85" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"61" , x"2A" , x"24" , x"24" , x"30" , x"80" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"68" , x"2F" , x"24" , x"25" , x"4F" , x"84" , x"5A" , x"2B" , x"24" , x"26" , x"4A" , x"87" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"84" , x"42" , x"25" , x"24" , x"24" , x"57" , x"8B" , x"92" , x"92" , x"92" , x"92" , x"92" , x"67" , x"2F" , x"24" , x"24" , x"24" , x"6D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7F" , x"3D" , x"24" , x"24" , x"24" , x"40" , x"32" , x"25" , x"24" , x"25" , x"36" , x"6E" , x"8E" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"73" , x"37" , x"25" , x"24" , x"2C" , x"65" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"70" , x"31" , x"25" , x"24" , x"33" , x"6C" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"78" , x"3D" , x"26" , x"24" , x"25" , x"4E" , x"87" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"58" , x"2B" , x"24" , x"24" , x"2E" , x"6C" , x"8E" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7D" , x"41" , x"26" , x"24" , x"24" , x"3F" , x"7B" , x"92" , x"92" , x"91" , x"57" , x"26" , x"24" , x"24" , x"3C" , x"83" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"90" , x"59" , x"2C" , x"24" , x"24" , x"37" , x"81" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"76" , x"31" , x"24" , x"24" , x"27" , x"6C" , x"8E" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8B" , x"56" , x"29" , x"24" , x"2B" , x"61" , x"8D" , x"74" , x"32" , x"24" , x"24" , x"38" , x"7B" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"74" , x"37" , x"24" , x"24" , x"2B" , x"6C" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"67" , x"2F" , x"24" , x"24" , x"24" , x"6D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7F" , x"3D" , x"24" , x"24" , x"24" , x"51" , x"55" , x"2E" , x"24" , x"24" , x"26" , x"46" , x"7C" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"73" , x"37" , x"25" , x"24" , x"2C" , x"65" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"6D" , x"31" , x"25" , x"24" , x"31" , x"6A" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"84" , x"4D" , x"31" , x"37" , x"38" , x"59" , x"88" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"58" , x"2B" , x"24" , x"24" , x"2E" , x"6C" , x"8E" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7E" , x"43" , x"26" , x"24" , x"24" , x"3C" , x"79" , x"92" , x"92" , x"8C" , x"50" , x"2B" , x"29" , x"26" , x"4B" , x"88" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"65" , x"2E" , x"24" , x"24" , x"32" , x"74" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8B" , x"3F" , x"26" , x"24" , x"25" , x"58" , x"89" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7D" , x"43" , x"25" , x"24" , x"37" , x"71" , x"90" , x"83" , x"42" , x"26" , x"24" , x"2E" , x"64" , x"8D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"63" , x"2E" , x"24" , x"24" , x"3A" , x"7A" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"67" , x"2F" , x"24" , x"24" , x"24" , x"6D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7F" , x"3D" , x"24" , x"24" , x"24" , x"54" , x"7C" , x"4F" , x"2A" , x"24" , x"24" , x"2A" , x"55" , x"87" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"73" , x"37" , x"25" , x"24" , x"2C" , x"65" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"73" , x"36" , x"25" , x"24" , x"27" , x"54" , x"88" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"90" , x"85" , x"80" , x"82" , x"82" , x"88" , x"90" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"58" , x"2B" , x"24" , x"24" , x"2E" , x"6C" , x"8E" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7C" , x"40" , x"26" , x"24" , x"24" , x"43" , x"7E" , x"92" , x"92" , x"8B" , x"70" , x"5F" , x"59" , x"52" , x"69" , x"8D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"61" , x"2D" , x"24" , x"24" , x"35" , x"7D" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"90" , x"4F" , x"29" , x"24" , x"25" , x"46" , x"85" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"6F" , x"34" , x"25" , x"25" , x"45" , x"81" , x"91" , x"88" , x"52" , x"2A" , x"24" , x"28" , x"56" , x"8A" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8A" , x"52" , x"28" , x"24" , x"24" , x"4C" , x"85" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"67" , x"2F" , x"24" , x"24" , x"24" , x"6D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7F" , x"3D" , x"24" , x"24" , x"24" , x"55" , x"8A" , x"75" , x"3C" , x"26" , x"24" , x"25" , x"32" , x"6B" , x"8F" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"73" , x"37" , x"25" , x"24" , x"2C" , x"65" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7E" , x"42" , x"26" , x"24" , x"25" , x"34" , x"65" , x"89" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"58" , x"2B" , x"24" , x"24" , x"2E" , x"6C" , x"8E" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"90" , x"71" , x"35" , x"25" , x"24" , x"24" , x"4E" , x"87" , x"92" , x"92" , x"91" , x"8E" , x"8D" , x"8C" , x"8A" , x"8D" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"4E" , x"29" , x"24" , x"25" , x"3D" , x"83" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"90" , x"62" , x"2D" , x"24" , x"24" , x"38" , x"7C" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8B" , x"5C" , x"2C" , x"24" , x"29" , x"55" , x"8A" , x"92" , x"8F" , x"66" , x"2E" , x"25" , x"25" , x"45" , x"80" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7F" , x"44" , x"26" , x"24" , x"2A" , x"5E" , x"8D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"67" , x"2F" , x"24" , x"24" , x"24" , x"6D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7F" , x"3D" , x"24" , x"24" , x"24" , x"55" , x"8B" , x"8B" , x"5F" , x"2E" , x"24" , x"24" , x"26" , x"40" , x"81" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"73" , x"37" , x"25" , x"24" , x"2C" , x"65" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8B" , x"58" , x"2A" , x"24" , x"24" , x"26" , x"35" , x"55" , x"6F" , x"87" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"58" , x"2B" , x"24" , x"24" , x"2E" , x"6C" , x"8E" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"87" , x"53" , x"2B" , x"24" , x"24" , x"2A" , x"5E" , x"8D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7C" , x"36" , x"25" , x"24" , x"25" , x"50" , x"87" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"7A" , x"37" , x"25" , x"24" , x"2F" , x"6B" , x"8E" , x"92" , x"92" , x"92" , x"92" , x"92" , x"85" , x"49" , x"28" , x"24" , x"30" , x"69" , x"8D" , x"92" , x"92" , x"78" , x"3B" , x"26" , x"24" , x"35" , x"6E" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"76" , x"39" , x"25" , x"24" , x"35" , x"6E" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"67" , x"2F" , x"24" , x"24" , x"24" , x"6D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7F" , x"3D" , x"24" , x"24" , x"24" , x"55" , x"8B" , x"91" , x"88" , x"4E" , x"28" , x"24" , x"24" , x"28" , x"56" , x"88" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"73" , x"37" , x"25" , x"24" , x"2C" , x"65" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"7E" , x"42" , x"25" , x"24" , x"24" , x"25" , x"28" , x"32" , x"3F" , x"54" , x"68" , x"7C" , x"88" , x"8C" , x"90" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"58" , x"2B" , x"24" , x"24" , x"2E" , x"6C" , x"8E" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"87" , x"5C" , x"31" , x"25" , x"24" , x"25" , x"3A" , x"74" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8A" , x"55" , x"29" , x"24" , x"24" , x"2C" , x"6F" , x"8E" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"85" , x"48" , x"28" , x"24" , x"2A" , x"5A" , x"8B" , x"92" , x"92" , x"92" , x"92" , x"91" , x"7C" , x"38" , x"26" , x"24" , x"39" , x"7B" , x"91" , x"92" , x"92" , x"84" , x"4B" , x"26" , x"24" , x"29" , x"5E" , x"8D" , x"92" , x"92" , x"92" , x"92" , x"91" , x"69" , x"2F" , x"24" , x"25" , x"42" , x"7D" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"67" , x"2F" , x"24" , x"24" , x"24" , x"6D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7F" , x"3D" , x"24" , x"24" , x"24" , x"55" , x"8B" , x"92" , x"92" , x"78" , x"3A" , x"25" , x"24" , x"25" , x"32" , x"68" , x"8C" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"73" , x"37" , x"25" , x"24" , x"2C" , x"65" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"90" , x"73" , x"3E" , x"28" , x"24" , x"24" , x"24" , x"24" , x"25" , x"29" , x"2E" , x"35" , x"41" , x"51" , x"65" , x"78" , x"80" , x"8A" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"58" , x"2B" , x"24" , x"24" , x"2E" , x"6C" , x"8E" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"84" , x"7B" , x"6F" , x"54" , x"2F" , x"25" , x"24" , x"24" , x"29" , x"56" , x"88" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8C" , x"67" , x"35" , x"25" , x"24" , x"24" , x"47" , x"85" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8A" , x"57" , x"2A" , x"24" , x"26" , x"4C" , x"87" , x"91" , x"92" , x"92" , x"92" , x"91" , x"66" , x"2F" , x"24" , x"26" , x"4D" , x"86" , x"92" , x"92" , x"92" , x"8E" , x"5B" , x"2A" , x"24" , x"25" , x"4C" , x"84" , x"92" , x"92" , x"92" , x"92" , x"8A" , x"55" , x"2A" , x"24" , x"27" , x"53" , x"89" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"67" , x"2F" , x"24" , x"24" , x"24" , x"6D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7F" , x"3D" , x"24" , x"24" , x"24" , x"55" , x"8B" , x"92" , x"92" , x"8D" , x"63" , x"31" , x"25" , x"24" , x"27" , x"42" , x"79" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"73" , x"37" , x"25" , x"24" , x"2C" , x"65" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8D" , x"72" , x"4A" , x"2D" , x"25" , x"24" , x"24" , x"24" , x"24" , x"24" , x"25" , x"26" , x"29" , x"2E" , x"37" , x"45" , x"56" , x"6D" , x"7F" , x"8F" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"58" , x"2B" , x"24" , x"24" , x"28" , x"43" , x"52" , x"54" , x"54" , x"54" , x"54" , x"54" , x"54" , x"54" , x"54" , x"54" , x"46" , x"3F" , x"34" , x"2A" , x"25" , x"24" , x"24" , x"25" , x"3E" , x"78" , x"8F" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8F" , x"70" , x"3D" , x"27" , x"24" , x"24" , x"32" , x"6C" , x"8F" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8F" , x"6A" , x"31" , x"25" , x"24" , x"3E" , x"7A" , x"90" , x"92" , x"92" , x"92" , x"90" , x"51" , x"29" , x"24" , x"26" , x"60" , x"8C" , x"92" , x"92" , x"92" , x"91" , x"6C" , x"32" , x"24" , x"24" , x"3A" , x"79" , x"92" , x"92" , x"92" , x"92" , x"84" , x"46" , x"27" , x"24" , x"2D" , x"62" , x"8D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"67" , x"2F" , x"24" , x"24" , x"24" , x"6D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7F" , x"3D" , x"24" , x"24" , x"24" , x"55" , x"8B" , x"92" , x"92" , x"92" , x"84" , x"4C" , x"28" , x"24" , x"24" , x"2A" , x"55" , x"88" , x"92" , x"92" , x"92" , x"92" , x"92" , x"73" , x"37" , x"25" , x"24" , x"2C" , x"65" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8E" , x"7F" , x"64" , x"41" , x"29" , x"25" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"25" , x"26" , x"29" , x"32" , x"43" , x"5F" , x"81" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"58" , x"2B" , x"24" , x"24" , x"24" , x"25" , x"25" , x"25" , x"25" , x"25" , x"25" , x"25" , x"25" , x"25" , x"25" , x"25" , x"25" , x"25" , x"24" , x"24" , x"24" , x"24" , x"27" , x"3D" , x"78" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8E" , x"6C" , x"3C" , x"27" , x"24" , x"25" , x"31" , x"61" , x"8B" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7B" , x"3F" , x"26" , x"24" , x"32" , x"6C" , x"90" , x"92" , x"92" , x"92" , x"85" , x"39" , x"24" , x"24" , x"2C" , x"7B" , x"91" , x"92" , x"92" , x"92" , x"92" , x"7F" , x"3E" , x"24" , x"24" , x"29" , x"6B" , x"91" , x"92" , x"92" , x"91" , x"7B" , x"35" , x"25" , x"24" , x"37" , x"79" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"67" , x"2F" , x"24" , x"24" , x"24" , x"6D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7F" , x"3D" , x"24" , x"24" , x"24" , x"55" , x"8B" , x"92" , x"92" , x"92" , x"91" , x"77" , x"3F" , x"27" , x"24" , x"24" , x"2E" , x"68" , x"8F" , x"92" , x"92" , x"92" , x"92" , x"73" , x"37" , x"25" , x"24" , x"2C" , x"65" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"8E" , x"85" , x"76" , x"58" , x"41" , x"32" , x"2C" , x"28" , x"25" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"25" , x"2B" , x"3E" , x"6A" , x"8A" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"58" , x"2B" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"27" , x"32" , x"4B" , x"76" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8A" , x"6D" , x"3A" , x"26" , x"24" , x"24" , x"2E" , x"56" , x"83" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"85" , x"4B" , x"26" , x"24" , x"2B" , x"61" , x"8E" , x"92" , x"92" , x"92" , x"6F" , x"2F" , x"24" , x"24" , x"3E" , x"85" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8F" , x"50" , x"26" , x"24" , x"25" , x"52" , x"8A" , x"92" , x"92" , x"90" , x"64" , x"2E" , x"24" , x"25" , x"46" , x"85" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"67" , x"2F" , x"24" , x"24" , x"24" , x"6D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7F" , x"3D" , x"24" , x"24" , x"24" , x"55" , x"8B" , x"92" , x"92" , x"92" , x"92" , x"8E" , x"67" , x"31" , x"24" , x"24" , x"25" , x"3D" , x"7C" , x"91" , x"92" , x"92" , x"92" , x"73" , x"37" , x"25" , x"24" , x"2C" , x"65" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"8A" , x"84" , x"75" , x"62" , x"52" , x"42" , x"35" , x"2C" , x"25" , x"24" , x"24" , x"24" , x"24" , x"24" , x"25" , x"35" , x"62" , x"87" , x"91" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"58" , x"2B" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"29" , x"2F" , x"37" , x"43" , x"57" , x"6C" , x"81" , x"8F" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8A" , x"64" , x"39" , x"25" , x"24" , x"24" , x"2A" , x"56" , x"81" , x"8F" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8E" , x"5E" , x"2B" , x"24" , x"25" , x"51" , x"88" , x"92" , x"92" , x"92" , x"5C" , x"29" , x"24" , x"24" , x"55" , x"8C" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"63" , x"2B" , x"24" , x"24" , x"3F" , x"85" , x"92" , x"92" , x"90" , x"51" , x"2A" , x"24" , x"26" , x"5A" , x"8A" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"67" , x"2F" , x"24" , x"24" , x"24" , x"6D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7F" , x"3D" , x"24" , x"24" , x"24" , x"55" , x"8B" , x"92" , x"92" , x"92" , x"92" , x"92" , x"86" , x"4F" , x"28" , x"24" , x"24" , x"29" , x"53" , x"86" , x"91" , x"92" , x"92" , x"73" , x"37" , x"25" , x"24" , x"2C" , x"65" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"90" , x"8D" , x"8A" , x"81" , x"71" , x"63" , x"53" , x"40" , x"2E" , x"24" , x"24" , x"24" , x"24" , x"26" , x"37" , x"6B" , x"8E" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"58" , x"2B" , x"24" , x"24" , x"2B" , x"51" , x"66" , x"68" , x"68" , x"68" , x"68" , x"68" , x"68" , x"68" , x"68" , x"68" , x"6B" , x"71" , x"76" , x"7F" , x"8C" , x"90" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"89" , x"5D" , x"35" , x"26" , x"24" , x"25" , x"2A" , x"52" , x"83" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"6F" , x"35" , x"24" , x"24" , x"40" , x"7D" , x"92" , x"92" , x"8B" , x"4A" , x"26" , x"24" , x"29" , x"6A" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"78" , x"32" , x"24" , x"24" , x"2C" , x"79" , x"91" , x"92" , x"8D" , x"3E" , x"25" , x"24" , x"2A" , x"73" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"67" , x"2F" , x"24" , x"24" , x"24" , x"6D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7F" , x"3D" , x"24" , x"24" , x"24" , x"55" , x"8B" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"7C" , x"3B" , x"25" , x"24" , x"25" , x"33" , x"68" , x"8E" , x"92" , x"92" , x"73" , x"37" , x"25" , x"24" , x"2C" , x"65" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"90" , x"8E" , x"8A" , x"7D" , x"6D" , x"4A" , x"2D" , x"26" , x"24" , x"24" , x"26" , x"44" , x"80" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"58" , x"2B" , x"24" , x"24" , x"2E" , x"6C" , x"8E" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"90" , x"7E" , x"4A" , x"2D" , x"25" , x"24" , x"25" , x"34" , x"62" , x"88" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"81" , x"40" , x"24" , x"24" , x"32" , x"74" , x"92" , x"92" , x"78" , x"3A" , x"24" , x"24" , x"38" , x"78" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8C" , x"40" , x"26" , x"24" , x"26" , x"63" , x"8C" , x"92" , x"78" , x"32" , x"24" , x"24" , x"3B" , x"83" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"67" , x"2F" , x"24" , x"24" , x"24" , x"6D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7F" , x"3D" , x"24" , x"24" , x"24" , x"55" , x"8B" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"90" , x"66" , x"32" , x"25" , x"24" , x"25" , x"3D" , x"75" , x"8F" , x"92" , x"73" , x"37" , x"25" , x"24" , x"2C" , x"65" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"87" , x"68" , x"3A" , x"26" , x"24" , x"24" , x"29" , x"69" , x"8F" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"58" , x"2B" , x"24" , x"24" , x"2E" , x"6C" , x"8E" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8D" , x"72" , x"45" , x"29" , x"25" , x"24" , x"25" , x"3A" , x"63" , x"88" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"90" , x"50" , x"26" , x"24" , x"28" , x"67" , x"90" , x"92" , x"68" , x"2F" , x"24" , x"25" , x"4C" , x"85" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"90" , x"55" , x"2B" , x"24" , x"25" , x"52" , x"88" , x"92" , x"67" , x"2C" , x"24" , x"24" , x"4E" , x"88" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"67" , x"2F" , x"24" , x"24" , x"24" , x"6D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7F" , x"3D" , x"24" , x"24" , x"24" , x"55" , x"8B" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"85" , x"55" , x"2C" , x"24" , x"24" , x"29" , x"4F" , x"85" , x"92" , x"73" , x"37" , x"25" , x"24" , x"2C" , x"65" , x"90" , x"92" , x"92" , x"92" , x"91" , x"85" , x"79" , x"75" , x"72" , x"78" , x"8D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"8A" , x"61" , x"2F" , x"24" , x"24" , x"25" , x"53" , x"8A" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"58" , x"2B" , x"24" , x"24" , x"2E" , x"6C" , x"8E" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8D" , x"68" , x"3D" , x"29" , x"24" , x"24" , x"25" , x"3C" , x"6F" , x"8B" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"64" , x"2B" , x"24" , x"24" , x"53" , x"8B" , x"8B" , x"55" , x"28" , x"24" , x"29" , x"5F" , x"8E" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"90" , x"69" , x"2E" , x"24" , x"25" , x"40" , x"84" , x"92" , x"55" , x"28" , x"24" , x"27" , x"65" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"67" , x"2F" , x"24" , x"24" , x"24" , x"6D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7F" , x"3D" , x"24" , x"24" , x"24" , x"55" , x"8B" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"79" , x"40" , x"25" , x"24" , x"24" , x"2F" , x"66" , x"8E" , x"73" , x"37" , x"25" , x"24" , x"2C" , x"65" , x"90" , x"92" , x"92" , x"92" , x"8F" , x"63" , x"3F" , x"38" , x"34" , x"45" , x"82" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"84" , x"3E" , x"24" , x"24" , x"24" , x"48" , x"87" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"58" , x"2B" , x"24" , x"24" , x"2E" , x"6C" , x"8E" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"8D" , x"5F" , x"36" , x"26" , x"24" , x"25" , x"2B" , x"46" , x"73" , x"8E" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"77" , x"31" , x"24" , x"24" , x"42" , x"86" , x"7F" , x"46" , x"26" , x"24" , x"34" , x"6D" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7D" , x"3B" , x"25" , x"24" , x"34" , x"75" , x"85" , x"46" , x"25" , x"24" , x"32" , x"75" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"67" , x"2F" , x"24" , x"24" , x"24" , x"6D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7F" , x"3D" , x"24" , x"24" , x"24" , x"55" , x"8B" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8D" , x"68" , x"32" , x"25" , x"24" , x"25" , x"3A" , x"7B" , x"71" , x"37" , x"25" , x"24" , x"2C" , x"65" , x"90" , x"92" , x"92" , x"92" , x"8E" , x"5B" , x"2C" , x"25" , x"25" , x"34" , x"71" , x"8F" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"4D" , x"26" , x"24" , x"24" , x"41" , x"84" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"58" , x"2B" , x"24" , x"24" , x"2E" , x"6C" , x"8E" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"84" , x"59" , x"2E" , x"24" , x"24" , x"24" , x"31" , x"57" , x"7F" , x"8F" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8B" , x"3E" , x"26" , x"24" , x"32" , x"7E" , x"75" , x"38" , x"25" , x"25" , x"43" , x"7F" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"87" , x"4F" , x"29" , x"24" , x"2D" , x"64" , x"70" , x"38" , x"24" , x"24" , x"46" , x"80" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"67" , x"2F" , x"24" , x"24" , x"24" , x"6D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7F" , x"3D" , x"24" , x"24" , x"24" , x"55" , x"8B" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8D" , x"55" , x"29" , x"24" , x"24" , x"26" , x"4E" , x"64" , x"35" , x"25" , x"24" , x"2C" , x"65" , x"90" , x"92" , x"92" , x"92" , x"91" , x"6A" , x"2F" , x"24" , x"24" , x"2B" , x"5B" , x"8A" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"90" , x"4A" , x"26" , x"24" , x"24" , x"48" , x"87" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"58" , x"2B" , x"24" , x"24" , x"2E" , x"6C" , x"8E" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"86" , x"58" , x"31" , x"25" , x"24" , x"24" , x"32" , x"61" , x"85" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"90" , x"52" , x"29" , x"24" , x"29" , x"6D" , x"64" , x"2E" , x"24" , x"28" , x"52" , x"89" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8E" , x"61" , x"2C" , x"24" , x"2A" , x"5A" , x"62" , x"2F" , x"24" , x"26" , x"57" , x"8A" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"67" , x"2F" , x"24" , x"24" , x"24" , x"6D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7F" , x"3D" , x"24" , x"24" , x"24" , x"55" , x"8B" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7C" , x"3D" , x"26" , x"24" , x"24" , x"30" , x"46" , x"31" , x"25" , x"24" , x"2C" , x"65" , x"90" , x"92" , x"92" , x"92" , x"92" , x"7C" , x"3A" , x"25" , x"24" , x"25" , x"3F" , x"78" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7F" , x"3D" , x"24" , x"24" , x"24" , x"51" , x"8A" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"58" , x"2B" , x"24" , x"24" , x"2E" , x"6C" , x"8E" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8B" , x"5F" , x"32" , x"26" , x"24" , x"25" , x"39" , x"65" , x"8A" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"90" , x"66" , x"2E" , x"24" , x"26" , x"55" , x"4D" , x"29" , x"24" , x"2E" , x"64" , x"8C" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"73" , x"37" , x"25" , x"26" , x"4B" , x"52" , x"29" , x"24" , x"2E" , x"67" , x"8F" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"67" , x"2F" , x"24" , x"24" , x"24" , x"6D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7F" , x"3D" , x"24" , x"24" , x"24" , x"55" , x"8B" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8F" , x"6A" , x"33" , x"25" , x"24" , x"26" , x"2C" , x"29" , x"24" , x"24" , x"2C" , x"65" , x"90" , x"92" , x"92" , x"92" , x"92" , x"88" , x"51" , x"28" , x"24" , x"24" , x"2B" , x"4F" , x"84" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8C" , x"60" , x"2F" , x"24" , x"24" , x"29" , x"69" , x"8F" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"58" , x"2B" , x"24" , x"24" , x"2E" , x"6C" , x"8E" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"90" , x"65" , x"34" , x"26" , x"24" , x"27" , x"3E" , x"70" , x"8C" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7C" , x"38" , x"25" , x"26" , x"41" , x"38" , x"26" , x"24" , x"35" , x"78" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7F" , x"46" , x"26" , x"24" , x"37" , x"3B" , x"26" , x"24" , x"3B" , x"77" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"67" , x"2F" , x"24" , x"24" , x"24" , x"6D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7F" , x"3D" , x"24" , x"24" , x"24" , x"55" , x"8B" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"88" , x"55" , x"2B" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"2C" , x"65" , x"90" , x"92" , x"92" , x"92" , x"92" , x"90" , x"72" , x"3A" , x"26" , x"24" , x"24" , x"2A" , x"4B" , x"79" , x"8B" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"90" , x"87" , x"61" , x"36" , x"26" , x"24" , x"25" , x"41" , x"7F" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"58" , x"2B" , x"24" , x"24" , x"2E" , x"6C" , x"8E" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7C" , x"3B" , x"25" , x"24" , x"24" , x"37" , x"6D" , x"8C" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"85" , x"48" , x"28" , x"25" , x"2E" , x"29" , x"25" , x"25" , x"49" , x"85" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8A" , x"55" , x"28" , x"24" , x"2C" , x"2D" , x"25" , x"26" , x"4D" , x"86" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"67" , x"2F" , x"24" , x"24" , x"24" , x"6D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7F" , x"3D" , x"24" , x"24" , x"24" , x"55" , x"8B" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"7C" , x"45" , x"27" , x"24" , x"24" , x"24" , x"24" , x"24" , x"2C" , x"65" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8A" , x"5E" , x"2E" , x"24" , x"24" , x"24" , x"29" , x"3A" , x"58" , x"73" , x"81" , x"88" , x"8F" , x"91" , x"91" , x"8D" , x"87" , x"80" , x"70" , x"4F" , x"31" , x"25" , x"24" , x"25" , x"33" , x"68" , x"8D" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"58" , x"2B" , x"24" , x"24" , x"2E" , x"6C" , x"8E" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8D" , x"5A" , x"29" , x"24" , x"24" , x"24" , x"3B" , x"5B" , x"63" , x"63" , x"63" , x"63" , x"63" , x"63" , x"63" , x"63" , x"63" , x"63" , x"63" , x"63" , x"63" , x"63" , x"69" , x"83" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8B" , x"5B" , x"2A" , x"24" , x"26" , x"25" , x"24" , x"25" , x"5E" , x"8B" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"68" , x"31" , x"24" , x"25" , x"25" , x"24" , x"2A" , x"5C" , x"8B" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"67" , x"2F" , x"24" , x"24" , x"24" , x"6D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7F" , x"3D" , x"24" , x"24" , x"24" , x"55" , x"8B" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"90" , x"6C" , x"34" , x"24" , x"24" , x"24" , x"24" , x"24" , x"2C" , x"65" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"83" , x"4F" , x"2A" , x"25" , x"24" , x"24" , x"26" , x"2B" , x"36" , x"45" , x"53" , x"5E" , x"63" , x"63" , x"5C" , x"4F" , x"43" , x"33" , x"28" , x"25" , x"24" , x"25" , x"2D" , x"57" , x"85" , x"91" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"58" , x"2B" , x"24" , x"24" , x"2E" , x"6C" , x"8E" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"79" , x"3D" , x"25" , x"24" , x"24" , x"24" , x"26" , x"29" , x"2A" , x"2A" , x"2A" , x"2A" , x"2A" , x"2A" , x"2A" , x"2A" , x"2A" , x"2A" , x"2A" , x"2A" , x"2A" , x"2A" , x"35" , x"70" , x"8E" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"90" , x"6D" , x"31" , x"25" , x"24" , x"24" , x"24" , x"28" , x"75" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"78" , x"3A" , x"24" , x"24" , x"24" , x"24" , x"31" , x"6E" , x"8E" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"67" , x"2F" , x"24" , x"24" , x"24" , x"6D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7F" , x"3D" , x"24" , x"24" , x"24" , x"55" , x"8B" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"89" , x"54" , x"28" , x"24" , x"24" , x"24" , x"24" , x"2C" , x"65" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"7E" , x"51" , x"2E" , x"25" , x"24" , x"24" , x"24" , x"25" , x"26" , x"29" , x"29" , x"2A" , x"2A" , x"29" , x"28" , x"26" , x"25" , x"24" , x"24" , x"24" , x"2C" , x"56" , x"81" , x"8F" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"58" , x"2B" , x"24" , x"24" , x"2E" , x"6C" , x"8E" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"65" , x"2E" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"30" , x"6E" , x"8E" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7B" , x"3F" , x"26" , x"24" , x"24" , x"24" , x"3B" , x"84" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8E" , x"4B" , x"25" , x"24" , x"24" , x"25" , x"40" , x"82" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"67" , x"2F" , x"24" , x"24" , x"24" , x"6D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7F" , x"3D" , x"24" , x"24" , x"24" , x"55" , x"8B" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"84" , x"44" , x"27" , x"24" , x"24" , x"24" , x"2C" , x"65" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"87" , x"69" , x"42" , x"2D" , x"26" , x"25" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"25" , x"2B" , x"3F" , x"6A" , x"88" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"58" , x"2B" , x"24" , x"24" , x"2E" , x"6C" , x"8E" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8C" , x"57" , x"28" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"24" , x"30" , x"6E" , x"8E" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"87" , x"50" , x"27" , x"24" , x"24" , x"24" , x"51" , x"8A" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"5E" , x"2A" , x"24" , x"24" , x"26" , x"53" , x"88" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"67" , x"2F" , x"24" , x"24" , x"24" , x"6D" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7F" , x"3D" , x"24" , x"24" , x"24" , x"55" , x"8B" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"6B" , x"35" , x"25" , x"24" , x"24" , x"2C" , x"65" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"8D" , x"7E" , x"66" , x"4C" , x"3C" , x"34" , x"2D" , x"28" , x"25" , x"24" , x"24" , x"26" , x"29" , x"2F" , x"38" , x"4B" , x"64" , x"7D" , x"8D" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"73" , x"5B" , x"57" , x"57" , x"5D" , x"7D" , x"8F" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"8D" , x"6F" , x"59" , x"57" , x"57" , x"57" , x"57" , x"57" , x"57" , x"57" , x"57" , x"57" , x"57" , x"57" , x"57" , x"57" , x"57" , x"57" , x"57" , x"57" , x"57" , x"57" , x"57" , x"5D" , x"7E" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"90" , x"74" , x"5A" , x"57" , x"57" , x"57" , x"76" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7B" , x"5C" , x"57" , x"57" , x"58" , x"76" , x"8E" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"7B" , x"5D" , x"57" , x"57" , x"57" , x"7E" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"87" , x"65" , x"57" , x"57" , x"57" , x"71" , x"8E" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"88" , x"6A" , x"59" , x"57" , x"57" , x"5C" , x"7B" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"90" , x"8E" , x"86" , x"78" , x"6E" , x"64" , x"5E" , x"58" , x"57" , x"57" , x"59" , x"5F" , x"67" , x"74" , x"86" , x"8D" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"90" , x"8D" , x"8E" , x"8E" , x"8D" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"8F" , x"8E" , x"8E" , x"8E" , x"8E" , x"8E" , x"8E" , x"8E" , x"8E" , x"8E" , x"8E" , x"8E" , x"8E" , x"8E" , x"8E" , x"8E" , x"8E" , x"8E" , x"8E" , x"8E" , x"8E" , x"8E" , x"8D" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"90" , x"8E" , x"8E" , x"8E" , x"8E" , x"90" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"8D" , x"8E" , x"8E" , x"8E" , x"90" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"8D" , x"8E" , x"8E" , x"8E" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"8E" , x"8E" , x"8E" , x"8E" , x"90" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"8F" , x"8E" , x"8E" , x"8E" , x"8E" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"91" , x"91" , x"90" , x"8E" , x"8E" , x"8E" , x"8E" , x"8E" , x"8E" , x"8E" , x"8F" , x"91" , x"91" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" ),
( x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" , x"92" )
);




END ImagePackage;

PACKAGE BODY ImagePackage IS

    
END PACKAGE BODY;